
`timescale 1ns/1ns
`define TIMESCALE

`include "sys_sig.v"

module fmul_top();

wire clk, reset;

sys_sig sys_sig (clk, reset);

reg [31:0] op1, op2;
reg [31:0] res_eth;

real op1_real, op2_real;
real res_eth_real;




FMUL32 #(.DATA_W(32), .OPERATION_NUM(4)) fmul
(
        .clk    (clk),
        .op1    (op1),
        .op2    (op2),
        .opc    (opcode),
        .r_mode (rmode),
        .result (result),
        .val    ()
);


always @(posedge clk) begin
op1 <= 32'b01100100001100010000010111101110;
op2 <= 32'b01010010111010010010001011010111;
#4;
op1 <= 32'b00010010010011010011001101011011;
op2 <= 32'b01000111111111011001010011011110;
#4;
op1 <= 32'b00111111101010011100111011001100;
op2 <= 32'b00111100011001100101000010110110;
#4;
op1 <= 32'b01101101111110110100011011101110;
op2 <= 32'b01110001110000011001011011010110;
#4;
op1 <= 32'b00011011111000010011100010100101;
op2 <= 32'b00100110100011010010010000100000;
#4;
op1 <= 32'b01001001101010010001010001111011;
op2 <= 32'b01011011001111001011010000001100;
#4;
op1 <= 32'b00110110110110100000101011110010;
op2 <= 32'b00001111100000101011100011110000;
#4;
op1 <= 32'b00100100110101111111011010000100;
op2 <= 32'b01000100100001011000001001101010;
#4;
op1 <= 32'b01010010100101010110010110001111;
op2 <= 32'b01111001000110110111010000101001;
#4;
op1 <= 32'b00000001011010011100010011000010;
op2 <= 32'b01101111001001010011000001111001;
#4;
op1 <= 32'b00101110001100000001100110001111;
op2 <= 32'b01100010110110101011101101010101;
#4;
op1 <= 32'b00011100011101010100000011010001;
op2 <= 32'b01011000001111111001011101001011;
#4;
op1 <= 32'b00001001110001110111000000111000;
op2 <= 32'b01001100011010110111111110100111;
#4;
op1 <= 32'b01111000101001100001101010110111;
op2 <= 32'b00000010001101101110101111011000;
#4;
op1 <= 32'b00100101100111001111001101111011;
op2 <= 32'b00110110011000110010001000000111;
#4;
op1 <= 32'b01010011101101000011000111101101;
op2 <= 32'b00101011010111100000000000100010;
#4;
op1 <= 32'b01000010000000000101101110000010;
op2 <= 32'b00100000101101010000000001000101;
#4;
op1 <= 32'b01101111101111100111001110101010;
op2 <= 32'b00010101011110011000110111110111;
#4;
op1 <= 32'b00011101101111000100100000010111;
op2 <= 32'b01001010100110000111000010010001;
#4;
op1 <= 32'b01001011100000111111001100100010;
op2 <= 32'b01111111000011001011100100011100;
#4;
op1 <= 32'b01111001001101110100001011100100;
op2 <= 32'b00110011110111011100101100110110;
#4;
op1 <= 32'b01100111011010011011111111010001;
op2 <= 32'b00101001000010101011101100111100;
#4;
op1 <= 32'b01010101011111101000101100001011;
op2 <= 32'b01011110001010001001000000101000;
#4;
op1 <= 32'b00000010101110001100101100000001;
op2 <= 32'b01010010010100001101101011110000;
#4;
op1 <= 32'b01110001000100101101000011101100;
op2 <= 32'b01000111111011010101000111101110;
#4;
op1 <= 32'b00011110101111111001100111100101;
op2 <= 32'b01111100011111011010110111000011;
#4;
op1 <= 32'b01001100110010011111010011111110;
op2 <= 32'b01110001110101101100110000100010;
#4;
op1 <= 32'b00111010001010101110010011100110;
op2 <= 32'b01100101111000100000111110111110;
#4;
op1 <= 32'b00101000110101111100111000010010;
op2 <= 32'b00011011100111110001111111100101;
#4;
op1 <= 32'b00010101110101000111110101001001;
op2 <= 32'b00001111100001110111111000001011;
#4;
op1 <= 32'b00000011011011110101010100001111;
op2 <= 32'b01000100001010100101110001101010;
#4;
op1 <= 32'b00110010001011110000100001001000;
op2 <= 32'b01111001111111001110001010010111;
#4;
op1 <= 32'b00011111111000000000100011110100;
op2 <= 32'b01101110100110000101010011001111;
#4;
op1 <= 32'b00001101111111001000010111100101;
op2 <= 32'b01100011101101110101110111101000;
#4;
op1 <= 32'b00111011100110000111001001110001;
op2 <= 32'b00011000011000010000111111010011;
#4;
op1 <= 32'b00101001001111011011000000111110;
op2 <= 32'b01001101000111011110111010000011;
#4;
op1 <= 32'b00010111010110000011100001100010;
op2 <= 32'b00000001110011011001011000110101;
#4;
op1 <= 32'b01000101110100001001111110010111;
op2 <= 32'b00110111100000111111001101010101;
#4;
op1 <= 32'b00110010101110011101000010000001;
op2 <= 32'b00101011011110110001101010111100;
#4;
op1 <= 32'b01100001010101000111011000000000;
op2 <= 32'b00100001001110001001101011101010;
#4;
op1 <= 32'b00001111010100110010111110101011;
op2 <= 32'b00010110000001100001101111010010;
#4;
op1 <= 32'b01111101000000001001110010011001;
op2 <= 32'b00001010100111001111100010101101;
#4;
op1 <= 32'b01101010011100010011010110011011;
op2 <= 32'b01111111001000101011011111110101;
#4;
op1 <= 32'b01011000001111000110100001110000;
op2 <= 32'b00110100000000101000010111110101;
#4;
op1 <= 32'b01000110001110111100111011000010;
op2 <= 32'b01101000111000101111010101001001;
#4;
op1 <= 32'b01110100010100110111000101001111;
op2 <= 32'b00011101111100001000111001000001;
#4;
op1 <= 32'b00100010010001110011001110010111;
op2 <= 32'b01010010111000001101001110010010;
#4;
op1 <= 32'b00001111111010101110000001010100;
op2 <= 32'b01000111101101001100010001101010;
#4;
op1 <= 32'b00111101110011110011101100000010;
op2 <= 32'b00111100100111010110110101000001;
#4;
op1 <= 32'b00101011101010101100101010101111;
op2 <= 32'b01110001010100110101010001110111;
#4;
op1 <= 32'b00011010010000010101100011100101;
op2 <= 32'b00100110111101111111100110111100;
#4;
op1 <= 32'b00000111000110110011001111100011;
op2 <= 32'b01011010101011110110001010111010;
#4;
op1 <= 32'b01110101100110110010111011001100;
op2 <= 32'b01010000011110011101110101010100;
#4;
op1 <= 32'b01100011001011001001010010010001;
op2 <= 32'b00000100111110000110011001110001;
#4;
op1 <= 32'b01010000110110001111110111000010;
op2 <= 32'b01111001010101011111110001110011;
#4;
op1 <= 32'b00111111000100101101011001001011;
op2 <= 32'b00101110111011000100000010110111;
#4;
op1 <= 32'b01101100101011000101000010010100;
op2 <= 32'b00100011100000000001101111010011;
#4;
op1 <= 32'b01011010101110010001011011010001;
op2 <= 32'b00011000011101011110000001110011;
#4;
op1 <= 32'b01001000100001010111101111101111;
op2 <= 32'b01001101010000101101101100101001;
#4;
op1 <= 32'b00110110100110011011111100000010;
op2 <= 32'b01000010010101100011110111000110;
#4;
op1 <= 32'b01100100010000110001111010010101;
op2 <= 32'b01110110111111010110010001110000;
#4;
op1 <= 32'b00010010011110000011000010011000;
op2 <= 32'b01101100001100000101111100100111;
#4;
op1 <= 32'b00000000010101011011011010000111;
op2 <= 32'b00100001000111110001111110011110;
#4;
op1 <= 32'b01101110001011010100001000100001;
op2 <= 32'b00010101111111110010111100101101;
#4;
op1 <= 32'b00011011110010100001001110010101;
op2 <= 32'b01001010100100011111000100001010;
#4;
op1 <= 32'b01001010010110001111010101001010;
op2 <= 32'b00000000001110000111100000100111;
#4;
op1 <= 32'b01110111101001000110001011001110;
op2 <= 32'b00110100001101010001010011100100;
#4;
op1 <= 32'b00100100111010000110011100101110;
op2 <= 32'b01101000101100010110111110000110;
#4;
op1 <= 32'b00010011101000000110111110010011;
op2 <= 32'b01011110011001100101100010000101;
#4;
op1 <= 32'b00000001001010100101100000100111;
op2 <= 32'b00010010101100111110111101010110;
#4;
op1 <= 32'b00101110111011010011001010110110;
op2 <= 32'b00000111110100101101011111010111;
#4;
op1 <= 32'b00011100101011111000001010111111;
op2 <= 32'b01111100100110101111101001011111;
#4;
op1 <= 32'b00001010011010000000100011010001;
op2 <= 32'b00110001000100011111101100010100;
#4;
op1 <= 32'b00111000100110001111111110100000;
op2 <= 32'b01100110010001110111111011110001;
#4;
op1 <= 32'b00100110011111011101111001011001;
op2 <= 32'b01011011001111000100111111111100;
#4;
op1 <= 32'b01010011111000001111111010000101;
op2 <= 32'b00001111100101001000010001001001;
#4;
op1 <= 32'b00000001111110100111010100101001;
op2 <= 32'b00000100110101100001001010000100;
#4;
op1 <= 32'b00110000010010111001110111110011;
op2 <= 32'b00111001111111000101011100010110;
#4;
op1 <= 32'b01011110010011001101001010000010;
op2 <= 32'b00101110111011101001001001110010;
#4;
op1 <= 32'b01001011110100011111101101000100;
op2 <= 32'b01100011101000000011101010011000;
#4;
op1 <= 32'b00111001101111101011000010101101;
op2 <= 32'b01011000011110001000110111001100;
#4;
op1 <= 32'b00101000000101111100110011101100;
op2 <= 32'b01001101111010101011010100110000;
#4;
op1 <= 32'b00010101101000011011001110100101;
op2 <= 32'b00000010010100011000101011000110;
#4;
op1 <= 32'b00000011100010011111000100011111;
op2 <= 32'b01110111011010010111010101000001;
#4;
op1 <= 32'b01110001000001010011111100100111;
op2 <= 32'b01101011110111101010100100000011;
#4;
op1 <= 32'b01011110110100101011100001010001;
op2 <= 32'b00100000101101101100000000000111;
#4;
op1 <= 32'b01001101101100011111101000111110;
op2 <= 32'b00010110100000110000111010010010;
#4;
op1 <= 32'b00111010111100000100101110000101;
op2 <= 32'b00001010110111000010010000010101;
#4;
op1 <= 32'b00101000010111100010101000111010;
op2 <= 32'b00111111001010011111010101001111;
#4;
op1 <= 32'b00010110011101110010111000101011;
op2 <= 32'b01110100011001000010101111011101;
#4;
op1 <= 32'b00000100011010010000010100111001;
op2 <= 32'b01101001000110110100101011011000;
#4;
op1 <= 32'b00110010001111010001111110001000;
op2 <= 32'b01011110000001000111110111011000;
#4;
op1 <= 32'b00011111111001111110100101101001;
op2 <= 32'b00010010101010111001101001010010;
#4;
op1 <= 32'b00001110000000100001100111000101;
op2 <= 32'b01000111111000011111011011110000;
#4;
op1 <= 32'b00111100001001001101100111011101;
op2 <= 32'b00111100110101010011001001001111;
#4;
op1 <= 32'b00101001111011010000100000001101;
op2 <= 32'b01110001100101011011111001010100;
#4;
op1 <= 32'b00010111110000110001001100011010;
op2 <= 32'b01100110011010011010010101000011;
#4;
op1 <= 32'b01000101100100011011111111110000;
op2 <= 32'b01011011001011000010001001001001;
#4;
op1 <= 32'b01110011011100010110111111100010;
op2 <= 32'b00010000001011110111101101001001;
#4;
op1 <= 32'b01100001000101011010011010010111;
op2 <= 32'b01000100111000111010101111010001;
#4;
op1 <= 32'b00001111010001111100110000011101;
op2 <= 32'b01111001111111100100111110010110;
#4;
op1 <= 32'b01111100101110000001000001010100;
op2 <= 32'b01101110101000011001100100000101;
#4;
op1 <= 32'b01101011000010001100110111111011;
op2 <= 32'b01100011110011010010010100010101;
#4;
op1 <= 32'b00011001010100010000111100110110;
op2 <= 32'b01011001000100000101010011100101;
#4;
op1 <= 32'b01000110011000110011000011101000;
op2 <= 32'b01001101001110011010010011000110;
#4;
op1 <= 32'b01110100111011010101100111101100;
op2 <= 32'b01000010101101100101010000001010;
#4;
op1 <= 32'b00100010011001001111100111000011;
op2 <= 32'b01110111001001100111010001110001;
#4;
op1 <= 32'b01010000001111011100110111010011;
op2 <= 32'b01101011111010000001000101011001;
#4;
op1 <= 32'b01111110000000010000101010011011;
op2 <= 32'b01100001000001110010001001011111;
#4;
op1 <= 32'b01101100100011010100111101000011;
op2 <= 32'b00010110001010100101101100101010;
#4;
op1 <= 32'b01011001111110010001001111101010;
op2 <= 32'b00001010111010111100010111111101;
#4;
op1 <= 32'b00001000001001101001110100011100;
op2 <= 32'b01111111111110110000100101000010;
#4;
op1 <= 32'b00110101100111011100110100011010;
op2 <= 32'b01110100100110100000111000011100;
#4;
op1 <= 32'b00100011101011010110101010010111;
op2 <= 32'b00101001011111000011110111101000;
#4;
op1 <= 32'b00010001011100001100000100001001;
op2 <= 32'b01011110001110000010001001000000;
#4;
op1 <= 32'b00111111100000111101011100110101;
op2 <= 32'b01010011010001010111000110011110;
#4;
op1 <= 32'b01101100101010101111100110100001;
op2 <= 32'b00000111101101100001101001110010;
#4;
op1 <= 32'b00011010110010000000000111100010;
op2 <= 32'b01111100101100011100101011100000;
#4;
op1 <= 32'b01001000110011010011101010111110;
op2 <= 32'b00110001101010011101000011110111;
#4;
op1 <= 32'b00110110101110001011010100011111;
op2 <= 32'b01100110001110011100011111100010;
#4;
op1 <= 32'b01100100011111111011111000101101;
op2 <= 32'b00011011011110010010101101110110;
#4;
op1 <= 32'b01010010010110101101010111110000;
op2 <= 32'b00010000001110100001011010010111;
#4;
op1 <= 32'b00000000010110100000010011101011;
op2 <= 32'b01000101000111011011100100111001;
#4;
op1 <= 32'b00101110100111001010101111101011;
op2 <= 32'b01111010100011111011010010100100;
#4;
op1 <= 32'b01011100000100101010110000001101;
op2 <= 32'b00101111000001001010011110110011;
#4;
op1 <= 32'b00001010001100110000011111111010;
op2 <= 32'b01100100000110101011110100001011;
#4;
op1 <= 32'b00110111100010000000011010100101;
op2 <= 32'b01011000010110000100001100011111;
#4;
op1 <= 32'b01100101111110101001111011010110;
op2 <= 32'b00001101101101110110101101000000;
#4;
op1 <= 32'b00010011011001010111101001011101;
op2 <= 32'b01000010001110110000011101100001;
#4;
op1 <= 32'b00000001000101010111011000111100;
op2 <= 32'b00110111000011111100101011101011;
#4;
op1 <= 32'b01101110111011001000110101110001;
op2 <= 32'b01101011101101001000011010110001;
#4;
op1 <= 32'b01011101010000111100000000001001;
op2 <= 32'b00100001001101011010010011110111;
#4;
op1 <= 32'b00001010111001100100110110010101;
op2 <= 32'b00010101101001001110110110010110;
#4;
op1 <= 32'b00111001000101010110110101111011;
op2 <= 32'b01001010111110111001010011100010;
#4;
op1 <= 32'b01100110111010110011110111011110;
op2 <= 32'b01111111100110111001101110011110;
#4;
op1 <= 32'b00010100010000011100001100000111;
op2 <= 32'b01110100000101010010001100001010;
#4;
op1 <= 32'b01000010110000111001011101101000;
op2 <= 32'b00101001011001010010001111101011;
#4;
op1 <= 32'b01110000011100101000101000000100;
op2 <= 32'b00011110001110110101001110110001;
#4;
op1 <= 32'b01011110101110111011101011010011;
op2 <= 32'b01010011110000110110001011000100;
#4;
op1 <= 32'b00001100000100110010111101101001;
op2 <= 32'b00000111111011100011101011001111;
#4;
op1 <= 32'b00111010100101011101010100010110;
op2 <= 32'b01111101011101001101101110111101;
#4;
op1 <= 32'b00100111101011101000111011010000;
op2 <= 32'b00110001100010011110011010011001;
#4;
op1 <= 32'b00010101100011111010100001100000;
op2 <= 32'b00100110011101000010101110101000;
#4;
op1 <= 32'b00000100000010010001000110000010;
op2 <= 32'b01011011111111001101101100011001;
#4;
op1 <= 32'b00110001101111101011111010001100;
op2 <= 32'b01010000101111111001001011001101;
#4;
op1 <= 32'b00011111000000001001000100011111;
op2 <= 32'b01000100110010111111001111110001;
#4;
op1 <= 32'b01001101110110111011010110110100;
op2 <= 32'b01111010111001100010001110011010;
#4;
op1 <= 32'b01111011000100100000010000110101;
op2 <= 32'b00101110111001101010010011101001;
#4;
op1 <= 32'b00101000111100101011100100001110;
op2 <= 32'b00100011110100111001111111100101;
#4;
op1 <= 32'b01010110011010000011100101010110;
op2 <= 32'b00011000011011000101010111000011;
#4;
op1 <= 32'b01000101000101000101101010000000;
op2 <= 32'b01001101110110101100101110001110;
#4;
op1 <= 32'b01110010101100111001110110011011;
op2 <= 32'b01000010011011111100001000010000;
#4;
op1 <= 32'b01100000101011011010010001101010;
op2 <= 32'b00110111011000110001010000100111;
#4;
op1 <= 32'b01001110010000100101001110000100;
op2 <= 32'b01101100001100011100011111000011;
#4;
op1 <= 32'b00111100000110110101111101000001;
op2 <= 32'b00100001000000011101000000110111;
#4;
op1 <= 32'b01101010100011100111011001100001;
op2 <= 32'b01010110010110101001100011011101;
#4;
op1 <= 32'b01011000000101111010000101010001;
op2 <= 32'b00001010101110010001110110100000;
#4;
op1 <= 32'b00000101111001111100101111011100;
op2 <= 32'b01111111110100110011011010001110;
#4;
op1 <= 32'b01110011011110001011110011000011;
op2 <= 32'b00110100010110100011100010110001;
#4;
op1 <= 32'b00100010000110111100110011011010;
op2 <= 32'b01101010000010001010111001110100;
#4;
op1 <= 32'b00001111011011110011010111101000;
op2 <= 32'b01011110001010000100001000010111;
#4;
op1 <= 32'b01111101001000000111011110110101;
op2 <= 32'b00010011000101110000100101001011;
#4;
op1 <= 32'b00101011001101010110000000001001;
op2 <= 32'b01001000001000001110011111101000;
#4;
op1 <= 32'b00011000101001101010000001000011;
op2 <= 32'b00111100011011111010101100111001;
#4;
op1 <= 32'b00000111101000100100100010101000;
op2 <= 32'b00110010010111001000010011100110;
#4;
op1 <= 32'b01110100110001001110001101111000;
op2 <= 32'b00100110101001010101110100100110;
#4;
op1 <= 32'b01100010001111111111111000110000;
op2 <= 32'b00011010111110111100011111101001;
#4;
op1 <= 32'b00010000101011100010101101111000;
op2 <= 32'b01010000100100111000001000011110;
#4;
op1 <= 32'b00111110111001110111111001110110;
op2 <= 32'b00000101110010000101010110010111;
#4;
op1 <= 32'b00101100101001011000010100001001;
op2 <= 32'b00111010011100011101110100000100;
#4;
op1 <= 32'b01011010101101100100001000101011;
op2 <= 32'b01101111101100111000010110001001;
#4;
op1 <= 32'b00001000001100000010001000000011;
op2 <= 32'b01100100000100101100101010011111;
#4;
op1 <= 32'b01110110011011011010010011011010;
op2 <= 32'b00011001010011001110000000100000;
#4;
op1 <= 32'b00100100000011010000110001110101;
op2 <= 32'b00001101111011011101001110111011;
#4;
op1 <= 32'b01010001111101011100011011000101;
op2 <= 32'b01000010111111010100011100011000;
#4;
op1 <= 32'b00111111111110111000100100100000;
op2 <= 32'b00110111110001100110011000101110;
#4;
op1 <= 32'b01101101011010110001010100010000;
op2 <= 32'b00101100011000001011000101101101;
#4;
op1 <= 32'b01011011100101101110111110101010;
op2 <= 32'b00100001100110011000110100100001;
#4;
op1 <= 32'b01001001000100010101111001101000;
op2 <= 32'b00010101111101110110110110101010;
#4;
op1 <= 32'b00110110111100111111100001000011;
op2 <= 32'b01001010101111010010100111010100;
#4;
op1 <= 32'b01100101001110110100000010110011;
op2 <= 32'b00000000000100100001111110001111;
#4;
op1 <= 32'b01010010111000100111010011101110;
op2 <= 32'b01110100100101011011110001000111;
#4;
op1 <= 32'b00000000010100111110001001110010;
op2 <= 32'b01101001000011100011100010100011;
#4;
op1 <= 32'b00101110101000111000000100111110;
op2 <= 32'b01011110100001100010000010001001;
#4;
op1 <= 32'b00011100100011111100000111010111;
op2 <= 32'b01010011010110001100000100010100;
#4;
op1 <= 32'b00001010011101000101101100101000;
op2 <= 32'b00001000011001011110100101010000;
#4;
op1 <= 32'b00111000011011011011110110110101;
op2 <= 32'b00111101011000111100100101101101;
#4;
op1 <= 32'b00100110001100111101110000010110;
op2 <= 32'b01110010000100111001001101001010;
#4;
op1 <= 32'b00010100010001010100010110111001;
op2 <= 32'b01100111000100101100000111001000;
#4;
op1 <= 32'b01000010000010101010111010111110;
op2 <= 32'b00011011111001010100111011111001;
#4;
op1 <= 32'b01110000000010001010101101111110;
op2 <= 32'b00010001000000101101010110011101;
#4;
op1 <= 32'b00011101010000001010100101111111;
op2 <= 32'b01000100111111101000011001100001;
#4;
op1 <= 32'b00001011110010010110000110100010;
op2 <= 32'b00111010100011110111111000100100;
#4;
op1 <= 32'b00111001101111101101010000100001;
op2 <= 32'b01101111101011110101100100110011;
#4;
op1 <= 32'b00100110101101110000111000101100;
op2 <= 32'b00100011101001001111001000101111;
#4;
op1 <= 32'b00010100011111101010111100101000;
op2 <= 32'b00011000011010010101001001011000;
#4;
op1 <= 32'b01000011011010010000100011000000;
op2 <= 32'b01001110010101000001000000110000;
#4;
op1 <= 32'b00110000110110001110110011010100;
op2 <= 32'b00000010100100010000000000100000;
#4;
op1 <= 32'b01011110111110101111001110001011;
op2 <= 32'b00111000000000000011111010001100;
#4;
op1 <= 32'b01001100100110001110011010100000;
op2 <= 32'b01101100101101001010100010001111;
#4;
op1 <= 32'b00111010011011000111100000110100;
op2 <= 32'b01100001001001011100101100011011;
#4;
op1 <= 32'b01101000010110010101010011001100;
op2 <= 32'b01010110010100100111101110000010;
#4;
op1 <= 32'b01010101111001011101110001110010;
op2 <= 32'b00001010111001101111001101010110;
#4;
op1 <= 32'b00000100000100101000011101110100;
op2 <= 32'b00000000000010101010100010100001;
#4;
op1 <= 32'b00110001101010011011001111111101;
op2 <= 32'b01110100101001010000010110001001;
#4;
op1 <= 32'b00100000000101100100101011001001;
op2 <= 32'b00101001111100111011100111100111;
#4;
op1 <= 32'b00001101011011101111110011010001;
op2 <= 32'b01011110010100001001000100100001;
#4;
op1 <= 32'b00111011101111100100100001001010;
op2 <= 32'b01010011101100101001011000001001;
#4;
op1 <= 32'b01101001011110001110100111000111;
op2 <= 32'b01001000011110100000000111110110;
#4;
op1 <= 32'b00010111111010110110111001000010;
op2 <= 32'b01111101100101011101000111010101;
#4;
op1 <= 32'b01000101000101011101111111011101;
op2 <= 32'b01110001111110001001001110000100;
#4;
op1 <= 32'b01110011010000011011010110000010;
op2 <= 32'b00100111001010011001011010110001;
#4;
op1 <= 32'b01100000111101001000100110100110;
op2 <= 32'b00011011110101010001001101001000;
#4;
op1 <= 32'b01001110100100110001001100010100;
op2 <= 32'b01010000011011011010000110001001;
#4;
op1 <= 32'b01111100101000011010011101110101;
op2 <= 32'b00000101101110000001000011010101;
#4;
op1 <= 32'b01101010110000111100101001001000;
op2 <= 32'b01111010101010010110111010000111;
#4;
op1 <= 32'b00011000010011010100100101110000;
op2 <= 32'b01101111001111111010001011101111;
#4;
op1 <= 32'b00000110100100111101011111110110;
op2 <= 32'b01100100011110010110111101000011;
#4;
op1 <= 32'b01110011110110001100000011001101;
op2 <= 32'b00011000111011110010011011010111;
#4;
op1 <= 32'b01100001110110001000111100001100;
op2 <= 32'b00001101110010110101110101001000;
#4;
op1 <= 32'b01001111111011010000010111001111;
op2 <= 32'b00000010111000000110101111000010;
#4;
op1 <= 32'b00111101101011110100010011010010;
op2 <= 32'b01110111011101110100110101001110;
#4;
op1 <= 32'b00101011000111100000110110100110;
op2 <= 32'b00101100001111010111010001100100;
#4;
op1 <= 32'b00011001011011110000011011110011;
op2 <= 32'b00100001011010001111011000010010;
#4;
op1 <= 32'b00000111001110000000111001101011;
op2 <= 32'b01010110000010011001100110011000;
#4;
op1 <= 32'b00110101010111011000100001101100;
op2 <= 32'b01001011001101000000100000111001;
#4;
op1 <= 32'b01100010101010100100101010110010;
op2 <= 32'b01111111011111110110011101010011;
#4;
op1 <= 32'b01010000111010100001100001100111;
op2 <= 32'b01110100110111000000100100011000;
#4;
op1 <= 32'b01111110111111001011101010010000;
op2 <= 32'b00101001111010001111101011000110;
#4;
op1 <= 32'b01101100111110001110010001111010;
op2 <= 32'b01011110110001010000100100111000;
#4;
op1 <= 32'b00011011000100100101011101100110;
op2 <= 32'b01010100000110011111011011010000;
#4;
op1 <= 32'b01001000011000111101011100000101;
op2 <= 32'b00001000010110110001000110010011;
#4;
op1 <= 32'b01110110110110000110111110010100;
op2 <= 32'b00111101110010101100011010001110;
#4;
op1 <= 32'b01100100101010101100100000100111;
op2 <= 32'b00110010101011111001001010000110;
#4;
op1 <= 32'b00010010100011101111110111101011;
op2 <= 32'b01100111010100100001110111100101;
#4;
op1 <= 32'b00111111101000000011011111011100;
op2 <= 32'b00011011101110101110011011111100;
#4;
op1 <= 32'b01101101110011000111100000101000;
op2 <= 32'b01010000101101110111111001001111;
#4;
op1 <= 32'b01011011111110011000000011011111;
op2 <= 32'b00000101110110011111000010001101;
#4;
op1 <= 32'b01001001110001011101010011011001;
op2 <= 32'b01111010101100111000110101000101;
#4;
op1 <= 32'b01110111000001111110011111110110;
op2 <= 32'b00101110111100110001111001101010;
#4;
op1 <= 32'b00100101100010111001001110100001;
op2 <= 32'b01100100101000000010001010000101;
#4;
op1 <= 32'b00010011000010011111101101110100;
op2 <= 32'b01011000110110011101010110010001;
#4;
op1 <= 32'b01000001001100101111100111000000;
op2 <= 32'b00001101111100111111101101101110;
#4;
op1 <= 32'b01101110110000011011011110100111;
op2 <= 32'b01000010110000111110100000101000;
#4;
op1 <= 32'b00011100011010011011110100000100;
op2 <= 32'b01110111010000001101101001100001;
#4;
op1 <= 32'b00001010110100110001111001101001;
op2 <= 32'b01101100111001000010100010110101;
#4;
op1 <= 32'b00111001000010000010011011000100;
op2 <= 32'b00100001110100011011100100000010;
#4;
op1 <= 32'b00100110001101101101100010110010;
op2 <= 32'b01010110001110101011000011001100;
#4;
op1 <= 32'b01010011110000110110100101011111;
op2 <= 32'b00001010100111101010110000000011;
#4;
op1 <= 32'b00000010001011011101011110011010;
op2 <= 32'b00000000001100100001100101110100;
#4;
op1 <= 32'b00110000101101010101110010100010;
op2 <= 32'b01110101011111011010001101110000;
#4;
op1 <= 32'b01011110000001000110101010000010;
op2 <= 32'b00101010000100101000110101111100;
#4;
op1 <= 32'b00001011111001101000000010110100;
op2 <= 32'b01011110111011001001111111100111;
#4;
op1 <= 32'b01111010000011001111110011111010;
op2 <= 32'b00010100000000100111110111001100;
#4;
op1 <= 32'b01100111011110111011111001000000;
op2 <= 32'b01001000100100111101000101001011;
#4;
op1 <= 32'b01010101010101101001000010100110;
op2 <= 32'b00111101010111010000000010011110;
#4;
op1 <= 32'b00000011011100010000011100110111;
op2 <= 32'b01110010010011010011111010011100;
#4;
op1 <= 32'b01110001001010010110001111100000;
op2 <= 32'b00100111001110110101100111011000;
#4;
op1 <= 32'b00011111010011101100011100111000;
op2 <= 32'b00011100010110001110111011111000;
#4;
op1 <= 32'b00001100001100011100110010010111;
op2 <= 32'b01010000001000111111110000010010;
#4;
op1 <= 32'b00111010101011001110001010111001;
op2 <= 32'b00000101110010011100011111010000;
#4;
op1 <= 32'b01101000100110010110011110001001;
op2 <= 32'b01111010100100111001101110000010;
#4;
op1 <= 32'b01010110101101111000001110100101;
op2 <= 32'b01101111101101010101001101001001;
#4;
op1 <= 32'b01000100010010001000110110110000;
op2 <= 32'b00100100010111011000100101011110;
#4;
op1 <= 32'b01110010101101111100000101010011;
op2 <= 32'b01011001110010010101011000011011;
#4;
op1 <= 32'b01011111111011100101110101011110;
op2 <= 32'b00001101101000001100011100111000;
#4;
op1 <= 32'b01001110001101001100001001111110;
op2 <= 32'b00000011010010010010111101111101;
#4;
op1 <= 32'b01111011011110101010011111100011;
op2 <= 32'b00110111011110011010100011100011;
#4;
op1 <= 32'b00101001100101001000001110101111;
op2 <= 32'b00101100101100000010111111101001;
#4;
op1 <= 32'b01010111100000111111010101010011;
op2 <= 32'b00100001100000101111111011010101;
#4;
op1 <= 32'b01000101100011000000110010000011;
op2 <= 32'b00010110011101011111011001110111;
#4;
op1 <= 32'b00110011110111100100111001000001;
op2 <= 32'b01001011110100110001101100000011;
#4;
op1 <= 32'b00100000100100111011000011101100;
op2 <= 32'b00111111101000001000010011011001;
#4;
op1 <= 32'b00001111000001011101110000010001;
op2 <= 32'b00110100110111010100000000001001;
#4;
op1 <= 32'b01111100111100000111111000111110;
op2 <= 32'b00101001111001110010011011001100;
#4;
op1 <= 32'b01101011001111100111110001100101;
op2 <= 32'b01011111010001011100111100011011;
#4;
op1 <= 32'b00011000011110011001010101011000;
op2 <= 32'b01010011100110110111110110100010;
#4;
op1 <= 32'b00000110101101100010100111101110;
op2 <= 32'b00001000110100011111011110101001;
#4;
op1 <= 32'b00110100010101111111111100101110;
op2 <= 32'b01111101010000001100111000010000;
#4;
op1 <= 32'b00100010110000101010110111001111;
op2 <= 32'b00110010110100000001100010000110;
#4;
op1 <= 32'b00001111101100110111110110011001;
op2 <= 32'b01100110110000000000110011011100;
#4;
op1 <= 32'b01111110001101011101111111000110;
op2 <= 32'b01011100001011110011100011100100;
#4;
op1 <= 32'b00101100000110000010001111011001;
op2 <= 32'b00010000110101100011111000100111;
#4;
op1 <= 32'b00011010010101010101111100011010;
op2 <= 32'b01000110011001101110011110110001;
#4;
op1 <= 32'b00000111111010000101011101010011;
op2 <= 32'b01111010111000010010010101101001;
#4;
op1 <= 32'b01110101010011111010010010100110;
op2 <= 32'b00101111010110111110001000100101;
#4;
op1 <= 32'b00100011000110011011110000110101;
op2 <= 32'b00100100001001101100001110011001;
#4;
op1 <= 32'b01010001011111111001100001111111;
op2 <= 32'b01011001010100000100001111010011;
#4;
op1 <= 32'b01111111000001111000010001110100;
op2 <= 32'b01001101111110110011111001111101;
#4;
op1 <= 32'b01101100100100100101111011001001;
op2 <= 32'b00000010100001101100011110110101;
#4;
op1 <= 32'b01011011010010001000101000111010;
op2 <= 32'b01111000011000010101110010111110;
#4;
op1 <= 32'b00001000101000000001001100101100;
op2 <= 32'b01101100100011100010000010001011;
#4;
op1 <= 32'b01110111001110000000111110110011;
op2 <= 32'b00100010010111010001011000011111;
#4;
op1 <= 32'b01100100110001011000101001001011;
op2 <= 32'b01010110110011001011111100010101;
#4;
op1 <= 32'b01010010111100111100011011110101;
op2 <= 32'b00001011111100110101100111001000;
#4;
op1 <= 32'b00000000010011111000101101010011;
op2 <= 32'b00000000011000000001001010000011;
#4;
op1 <= 32'b00101110100010010011001010000010;
op2 <= 32'b01110101100100100100000111001100;
#4;
op1 <= 32'b01011100000111010100001100011000;
op2 <= 32'b01101010000101010100110010010010;
#4;
op1 <= 32'b01001010000001111010011100110010;
op2 <= 32'b01011111001000000011000001010001;
#4;
op1 <= 32'b01110111110001010101011010101010;
op2 <= 32'b00010011110000011011001110010101;
#4;
op1 <= 32'b00100101010110110111010000101101;
op2 <= 32'b00001000011110111110011111111001;
#4;
op1 <= 32'b01010011010111001101111011000011;
op2 <= 32'b00111101010011001000010000001010;
#4;
op1 <= 32'b01000001100011000101101101101100;
op2 <= 32'b00110010011100101001001011000000;
#4;
op1 <= 32'b00101111010001010011100111101110;
op2 <= 32'b00100111000010001110100111100000;
#4;
op1 <= 32'b00011100110010010101111011100010;
op2 <= 32'b01011011101100100111000000110100;
#4;
op1 <= 32'b01001011011100011111100100011110;
op2 <= 32'b00010001100010110000010100011100;
#4;
op1 <= 32'b00111001001011000011001001010101;
op2 <= 32'b01000110000000000100100111101001;
#4;
op1 <= 32'b00100111000010111111101101011110;
op2 <= 32'b00111011001001011111101111111010;
#4;
op1 <= 32'b00010100100110001101001011111001;
op2 <= 32'b00101111101111010001101101011111;
#4;
op1 <= 32'b01000010011001000101011011111000;
op2 <= 32'b00100100010100011110011110101001;
#4;
op1 <= 32'b01110000100101011010101100000100;
op2 <= 32'b00011001100010101001100011000111;
#4;
op1 <= 32'b00011110100011100110001010011010;
op2 <= 32'b01001110011100001111100011101110;
#4;
op1 <= 32'b00001100001000110001001110000011;
op2 <= 32'b00000010111101000110111100110000;
#4;
op1 <= 32'b00111010011000111010011111001111;
op2 <= 32'b00111000101001001110101010001000;
#4;
op1 <= 32'b00101000010001001101100000001100;
op2 <= 32'b01101101010101010011111000111111;
#4;
op1 <= 32'b00010110000000001011010101101110;
op2 <= 32'b01100001110111011011101101111110;
#4;
op1 <= 32'b01000011110010111011000111111101;
op2 <= 32'b00010110101111101101010011110111;
#4;
op1 <= 32'b01110001101000100100011110111010;
op2 <= 32'b00001011101111111011010010101001;
#4;
op1 <= 32'b00011111001101000100110111000111;
op2 <= 32'b01000000001101111010001110011100;
#4;
op1 <= 32'b00001101011001000010000000010011;
op2 <= 32'b01110101010001100011100010000011;
#4;
op1 <= 32'b01111011001110001110001110101011;
op2 <= 32'b01101010000101010011001101100100;
#4;
op1 <= 32'b00101001010100101110101110101000;
op2 <= 32'b01011111011010011010101110100001;
#4;
op1 <= 32'b01010110110011111111111001111011;
op2 <= 32'b01010011111101101101011011011001;
#4;
op1 <= 32'b00000101010101111000010001011000;
op2 <= 32'b01001001011111011001010010100110;
#4;
op1 <= 32'b00110011010000110111110011010011;
op2 <= 32'b01111110011001011001000101110011;
#4;
op1 <= 32'b01100000010011001000010100001010;
op2 <= 32'b00110010010100011111001111011010;
#4;
op1 <= 32'b01001110011100011010111010100000;
op2 <= 32'b00100111100111010101111011001010;
#4;
op1 <= 32'b00111100011110011101100000100000;
op2 <= 32'b01011100100001011010101001100000;
#4;
op1 <= 32'b00101010010110011011001001011001;
op2 <= 32'b00010001010010101010110100000011;
#4;
op1 <= 32'b00010111111011000101110100010011;
op2 <= 32'b00000110000011001010101100100101;
#4;
op1 <= 32'b00000101110010011101011010110111;
op2 <= 32'b01111010111011101100010010001010;
#4;
op1 <= 32'b01110011100110011110100100001001;
op2 <= 32'b01101111100011000111001110010101;
#4;
op1 <= 32'b01100001010000010001000101110100;
op2 <= 32'b00100100010110100001010001000101;
#4;
op1 <= 32'b00001110111001001011111101110100;
op2 <= 32'b00011000110011110000010000010001;
#4;
op1 <= 32'b01111101000100110011011000101100;
op2 <= 32'b01001110000001111011100101010010;
#4;
op1 <= 32'b00101010111110110111000000001111;
op2 <= 32'b01000011000000100010101110000111;
#4;
op1 <= 32'b00011001101011010000111000111100;
op2 <= 32'b01111000110011101100100111110110;
#4;
op1 <= 32'b01000111001011010110001110010000;
op2 <= 32'b00101101001011000100111010101111;
#4;
op1 <= 32'b00110101000010001010110001101101;
op2 <= 32'b00100010000100011000001100101100;
#4;
op1 <= 32'b00100011010110001111001110100111;
op2 <= 32'b00010111011100010010101101100000;
#4;
op1 <= 32'b01010001000011101101111001000001;
op2 <= 32'b00001011111010100010000111000001;
#4;
op1 <= 32'b00111110010010110011101011011011;
op2 <= 32'b01000000011111101010110111011000;
#4;
op1 <= 32'b00101100111000010010010101111011;
op2 <= 32'b01110101111101000110100000110000;
#4;
op1 <= 32'b01011010010100111101001101010101;
op2 <= 32'b01101010010001111101111110111111;
#4;
op1 <= 32'b00000111111111101000100111101000;
op2 <= 32'b01011111000100000100001001100111;
#4;
op1 <= 32'b01110101110000001101000110111011;
op2 <= 32'b00010100000010001101010010100001;
#4;
op1 <= 32'b01100011101101010101011110111100;
op2 <= 32'b01001000011111111001000100101000;
#4;
op1 <= 32'b01010001110111011100000000101011;
op2 <= 32'b01111110000000010111000001110110;
#4;
op1 <= 32'b01111111010011100010110111111000;
op2 <= 32'b01110010001111000101000100000001;
#4;
op1 <= 32'b00101101100000100111100101011011;
op2 <= 32'b01100111101011111011100010010101;
#4;
op1 <= 32'b00011010101000110110110111100111;
op2 <= 32'b00011011110010000001100011001101;
#4;
op1 <= 32'b01001001011010011111111010110001;
op2 <= 32'b00010001100010010000001101001111;
#4;
op1 <= 32'b01110111011110011100011100100110;
op2 <= 32'b00000110101000100110100010101010;
#4;
op1 <= 32'b00100100100100010110010011110011;
op2 <= 32'b01111010110111011110100011010110;
#4;
op1 <= 32'b01010010011001111001101111101011;
op2 <= 32'b01101111100110010001110011100010;
#4;
op1 <= 32'b01000000100000101010010011101110;
op2 <= 32'b00100100101110100010001111111010;
#4;
op1 <= 32'b00101111001110010101111101011010;
op2 <= 32'b00011010000110111000011111110110;
#4;
op1 <= 32'b00011100101101100100110011001000;
op2 <= 32'b01001110101111111011000010010001;
#4;
op1 <= 32'b00001010100101000100010001000000;
op2 <= 32'b00000011101010010101100101000011;
#4;
op1 <= 32'b01111000000110010110000000001011;
op2 <= 32'b00111000001001101110000111111001;
#4;
op1 <= 32'b01100110011111001100001110000000;
op2 <= 32'b01101101100110111110101101011100;
#4;
op1 <= 32'b01010100001000011100010111100011;
op2 <= 32'b01100001111110100001001100100110;
#4;
op1 <= 32'b01000001111011110000110011111010;
op2 <= 32'b00010110111010000010011001111011;
#4;
op1 <= 32'b00101111011001011111000010010000;
op2 <= 32'b00001011011001100110110001100111;
#4;
op1 <= 32'b00011101011111001101010100100100;
op2 <= 32'b01000000100011101011011011001001;
#4;
op1 <= 32'b00001011110011010100011110100111;
op2 <= 32'b01110101101001001000001100101111;
#4;
op1 <= 32'b01111001001111001011001111001110;
op2 <= 32'b01101010011011110001001010101000;
#4;
op1 <= 32'b01100111000010100100110010010010;
op2 <= 32'b00011111001010011010111110101001;
#4;
op1 <= 32'b00010100111110110110010000101101;
op2 <= 32'b00010011111111010111111011001011;
#4;
op1 <= 32'b01000011001111001111101110110110;
op2 <= 32'b01001001001111001011111100011001;
#4;
op1 <= 32'b01110000110010111110101011100010;
op2 <= 32'b01111101111110011101111000010101;
#4;
op1 <= 32'b01011111000100011100000011011110;
op2 <= 32'b00110011001000011111110101001010;
#4;
op1 <= 32'b00001011110110111010110011011110;
op2 <= 32'b00100110111110101110111000010011;
#4;
op1 <= 32'b01111010100001000011100011101100;
op2 <= 32'b00011100101000101011000000011010;
#4;
op1 <= 32'b01101000001010000000010001111110;
op2 <= 32'b00010001010010110000101100110111;
#4;
op1 <= 32'b01010110000111000111011000001011;
op2 <= 32'b00000110001100010010011101000100;
#4;
op1 <= 32'b00000011101010110011001111111000;
op2 <= 32'b00111010101111110000111110000110;
#4;
op1 <= 32'b01110010011000000100101010011011;
op2 <= 32'b00110000011110011100010111111101;
#4;
op1 <= 32'b00011111010110010110110011001000;
op2 <= 32'b01100100100000001110110000011111;
#4;
op1 <= 32'b00001101110011110111100010110011;
op2 <= 32'b00011001111110010101000000010000;
#4;
op1 <= 32'b01111011011011110111111011000100;
op2 <= 32'b01001110011000101001000010011011;
#4;
op1 <= 32'b01101001011000010000110000001010;
op2 <= 32'b00000011011001111010110010001110;
#4;
op1 <= 32'b00010111001010011110010101110101;
op2 <= 32'b01111000011111111011101100010111;
#4;
op1 <= 32'b00000101101001011110100011101110;
op2 <= 32'b01101101110101011010011000100110;
#4;
op1 <= 32'b00110011001100001010110001000001;
op2 <= 32'b01100010010110000101001111010110;
#4;
op1 <= 32'b00100000101101111110000110110001;
op2 <= 32'b01010110101111010100010011100101;
#4;
op1 <= 32'b00001110110101110111110110010111;
op2 <= 32'b00001100001010011011010101011101;
#4;
op1 <= 32'b01111100010111110001011110010011;
op2 <= 32'b01000000011100101011010100101011;
#4;
op1 <= 32'b01101010100101001000001111011101;
op2 <= 32'b01110101100100100001101000111001;
#4;
op1 <= 32'b01011000100100100001110111010111;
op2 <= 32'b00101010101101111100000101101010;
#4;
op1 <= 32'b01000110000000010001110001000011;
op2 <= 32'b01011111001001011011000010101010;
#4;
op1 <= 32'b00110011100000000101100101001111;
op2 <= 32'b00010011101111100110000010110101;
#4;
op1 <= 32'b00100001111011100001110100001100;
op2 <= 32'b00001000111000101101101100101011;
#4;
op1 <= 32'b00001111100011110001100010111000;
op2 <= 32'b01111101011100010101110100001010;
#4;
op1 <= 32'b01111101010110010111001100000001;
op2 <= 32'b01110010010100010011001101110001;
#4;
op1 <= 32'b01101011001100000100010111000111;
op2 <= 32'b01100111001011001100001010000000;
#4;
op1 <= 32'b01011001000100000011011101111011;
op2 <= 32'b00011100000010011001010000010011;
#4;
op1 <= 32'b01000111100000011011110010111100;
op2 <= 32'b01010001100110111001011011111001;
#4;
op1 <= 32'b00110101010010010000111011111001;
op2 <= 32'b00000110011111111010001011100001;
#4;
op1 <= 32'b01100011011101010101100110010000;
op2 <= 32'b00111011110000100101001001001111;
#4;
op1 <= 32'b00010001001010100100000100000101;
op2 <= 32'b01110000011011000000001010110101;
#4;
op1 <= 32'b01111111000011001000110111101101;
op2 <= 32'b01100101001011111100011101001001;
#4;
op1 <= 32'b01101100111111101001000111010000;
op2 <= 32'b01011001111111010101101100001000;
#4;
op1 <= 32'b00011010011011001100110011111010;
op2 <= 32'b01001110110010010111011111001111;
#4;
op1 <= 32'b00001000101010001101010000101111;
op2 <= 32'b00000011111101010100110011110111;
#4;
op1 <= 32'b00110110100000000100000110111100;
op2 <= 32'b01111000110011011101100100000010;
#4;
op1 <= 32'b00100100010110111000101100001001;
op2 <= 32'b00101101011001000100010111100000;
#4;
op1 <= 32'b00010001100111001100111001110110;
op2 <= 32'b00100001110101101000010011101101;
#4;
op1 <= 32'b00111111110010000111001010101010;
op2 <= 32'b00010110111111010111010001111111;
#4;
op1 <= 32'b00101101101011100000000011011110;
op2 <= 32'b00001011110011000111110111100110;
#4;
op1 <= 32'b01011011100100110110010001000110;
op2 <= 32'b00000000100111011010011000100001;
#4;
op1 <= 32'b00001001000111101011101100000100;
op2 <= 32'b01110101001101101000000000001010;
#4;
op1 <= 32'b01111000000110011100100001110101;
op2 <= 32'b01101011010110101000001100001011;
#4;
op1 <= 32'b00100101011000110111110110010000;
op2 <= 32'b00011111100001100010111101010100;
#4;
op1 <= 32'b00010011011001100010111001111010;
op2 <= 32'b01010100100110001000000111100000;
#4;
op1 <= 32'b01000001001010000101111101011000;
op2 <= 32'b00001001010000000100101100001110;
#4;
op1 <= 32'b01101110110101101000010000010001;
op2 <= 32'b01111110000000101100000101100111;
#4;
op1 <= 32'b01011100111110011100011000010100;
op2 <= 32'b01110011000111011110110100000011;
#4;
op1 <= 32'b01001010100111100111001111010001;
op2 <= 32'b01100111100110110001111111111111;
#4;
op1 <= 32'b01111000000111000110001010101100;
op2 <= 32'b00011100000101110001110000101100;
#4;
op1 <= 32'b00100110100101001010100100110000;
op2 <= 32'b01010001111000101100101101101001;
#4;
op1 <= 32'b00010100101001100100100010110001;
op2 <= 32'b00000110100111010101100100010110;
#4;
op1 <= 32'b00000010000111110100100110011101;
op2 <= 32'b01111011001011101110111010101110;
#4;
op1 <= 32'b01101111111101100000000011010100;
op2 <= 32'b01110000001000000110010001111100;
#4;
op1 <= 32'b01011110000001001001000000100010;
op2 <= 32'b00100100111100111000101000111101;
#4;
op1 <= 32'b00001011110000000010011101100010;
op2 <= 32'b01011001110010101011001001000101;
#4;
op1 <= 32'b01111001100011101001000100101010;
op2 <= 32'b01001110100001101101110110101011;
#4;
op1 <= 32'b01100111101101000011010011111101;
op2 <= 32'b01000011111111111100101011100000;
#4;
op1 <= 32'b01010101010001100011100000111110;
op2 <= 32'b00111000100110110011001110001100;
#4;
op1 <= 32'b00000011011100101101000000011000;
op2 <= 32'b00101101101010100111000111010100;
#4;
op1 <= 32'b00110001100001111110110010010110;
op2 <= 32'b01100010101111011000000100000010;
#4;
op1 <= 32'b00011110101001111100000000000011;
op2 <= 32'b00010110111000001111000010110000;
#4;
op1 <= 32'b01001100101010110111101110111101;
op2 <= 32'b00001011111001010110001101011100;
#4;
op1 <= 32'b01111011000110011101110111100110;
op2 <= 32'b00000001001110110111110100101011;
#4;
op1 <= 32'b01101000110001011110100100011000;
op2 <= 32'b00110101110110001111010010011011;
#4;
op1 <= 32'b01010110100101101011001000000000;
op2 <= 32'b00101010110001110000001111010000;
#4;
op1 <= 32'b00000100010101001011101011111000;
op2 <= 32'b01011111101010000000010000100110;
#4;
op1 <= 32'b01110001110101101001111101110001;
op2 <= 32'b01010011111011110111100111010011;
#4;
op1 <= 32'b01100000100010011010111011100100;
op2 <= 32'b00001001100010100010111101100011;
#4;
op1 <= 32'b01001101110011010110011111100010;
op2 <= 32'b01111110000010110001100111100100;
#4;
op1 <= 32'b01111011101100001100111000100000;
op2 <= 32'b01110010100101000111000010111001;
#4;
op1 <= 32'b01101001110010011100111010011100;
op2 <= 32'b00100111111011110001010111110110;
#4;
op1 <= 32'b01011000010100111101000111011100;
op2 <= 32'b01011101100101111010000010101000;
#4;
op1 <= 32'b01000101101100010010110101110000;
op2 <= 32'b00010001111000011010010111111100;
#4;
op1 <= 32'b01110011011000100111110100111001;
op2 <= 32'b00000110101101111100111100011011;
#4;
op1 <= 32'b00100001010111000111010111101010;
op2 <= 32'b00111011100100110101010001000110;
#4;
op1 <= 32'b00001111010011101011000101010000;
op2 <= 32'b01110000011101100100100010001001;
#4;
op1 <= 32'b01111101011111111110000101011000;
op2 <= 32'b00100101100011101001010110001111;
#4;
op1 <= 32'b01101010110011111110000011010110;
op2 <= 32'b01011001111110111110001011001000;
#4;
op1 <= 32'b01011000100111110111011001111001;
op2 <= 32'b01001110101011001101010100001100;
#4;
op1 <= 32'b01000110101101011010011101110101;
op2 <= 32'b01000011110101110100001111011001;
#4;
op1 <= 32'b00110101010011110100101100111001;
op2 <= 32'b00111001011011110011111111101100;
#4;
op1 <= 32'b01100010010100001101011111111101;
op2 <= 32'b00101101010101111111010000101001;
#4;
op1 <= 32'b01001111101110110100010101101001;
op2 <= 32'b01100001101110101101110000111110;
#4;
op1 <= 32'b01111110001111101010110001110011;
op2 <= 32'b01010111011001100000011100001011;
#4;
op1 <= 32'b01101011010000001010001101010010;
op2 <= 32'b01001011000110011101001110111110;
#4;
op1 <= 32'b01011001101011110111010101100111;
op2 <= 32'b00000000110011001110110011100000;
#4;
op1 <= 32'b01000111101101011001001100111001;
op2 <= 32'b00110101111101011011011110110110;
#4;
op1 <= 32'b00110101111011010001011011111110;
op2 <= 32'b00101011001011001011011001100000;
#4;
op1 <= 32'b01100011100001100100100011000011;
op2 <= 32'b01011111111010000001011010101111;
#4;
op1 <= 32'b01010001010010100101010010100001;
op2 <= 32'b00010100101000011111100000100111;
#4;
op1 <= 32'b00111111000000001011110011101010;
op2 <= 32'b00001001010000001111110010011101;
#4;
op1 <= 32'b00101101011010111011110110001100;
op2 <= 32'b01111110100010011000100001101101;
#4;
op1 <= 32'b01011011001101001001011001001111;
op2 <= 32'b00110011011100100101001000101010;
#4;
op1 <= 32'b01001001001000111110000001000000;
op2 <= 32'b00101000011101001110101001110101;
#4;
op1 <= 32'b00110111001011101001111110010000;
op2 <= 32'b01011101010110110000010100011110;
#4;
op1 <= 32'b00100100110001110000000010001000;
op2 <= 32'b00010001111100011110100101110000;
#4;
op1 <= 32'b00010010101110011101000011110011;
op2 <= 32'b01000110111000001001110101011100;
#4;
op1 <= 32'b01111111110110010101111110110011;
op2 <= 32'b01111010111100100100011100101010;
#4;
op1 <= 32'b00101110010000100101001000110000;
op2 <= 32'b01110000100100101001101111111000;
#4;
op1 <= 32'b00011100000110110110100101101100;
op2 <= 32'b00100101000010010011111101110010;
#4;
op1 <= 32'b00001010001100011101110100100100;
op2 <= 32'b01011010001000001000001100101010;
#4;
op1 <= 32'b01110111100010000100100001010110;
op2 <= 32'b00001110110110111100011100001111;
#4;
op1 <= 32'b01100110000110010101111100011001;
op2 <= 32'b01000100011101001101100001110101;
#4;
op1 <= 32'b01010011100000110101011100101100;
op2 <= 32'b01111000100111101111010111001111;
#4;
op1 <= 32'b00000001110101011101011001000001;
op2 <= 32'b01101110000011010110011001011110;
#4;
op1 <= 32'b01101111010001100000010010001010;
op2 <= 32'b01100010101010110100100001110001;
#4;
op1 <= 32'b00011100111010000100110001111110;
op2 <= 32'b01010110111110111111110101111100;
#4;
op1 <= 32'b00001010110001100011010101110011;
op2 <= 32'b00001100000101000111001100110111;
#4;
op1 <= 32'b01111000111000011011000011000010;
op2 <= 32'b00000000110100000001100111011111;
#4;
op1 <= 32'b01100110101101011110111010110111;
op2 <= 32'b00110110000001101001011000000111;
#4;
op1 <= 32'b01010100010101010110011101101010;
op2 <= 32'b00101010100010101110010001101101;
#4;
op1 <= 32'b01000010010000101111001101001100;
op2 <= 32'b00011111101000101111010000111001;
#4;
op1 <= 32'b01110000101011101100100111111100;
op2 <= 32'b01010100100110101011010001100110;
#4;
op1 <= 32'b00011101101100110101110001011000;
op2 <= 32'b01001000111100110100010010101011;
#4;
op1 <= 32'b01001011111110110110010100001010;
op2 <= 32'b01111110001010100101100001010000;
#4;
op1 <= 32'b00111010000010111100111010011110;
op2 <= 32'b00110011011000000111010100000000;
#4;
op1 <= 32'b01100111101000000111010100101010;
op2 <= 32'b00100111111011001110011010000010;
#4;
op1 <= 32'b01010110000110000100101010111001;
op2 <= 32'b01011101101000001000011101010010;
#4;
op1 <= 32'b00000011111110110111101001010110;
op2 <= 32'b00010010010010110111001110101001;
#4;
op1 <= 32'b00110001111010000100011110010111;
op2 <= 32'b01000111000101010110001101011111;
#4;
op1 <= 32'b01011111100100100111110010000110;
op2 <= 32'b00111011111100010010011010011000;
#4;
op1 <= 32'b00001101011000010111011011001100;
op2 <= 32'b00110000100001001110011010000110;
#4;
op1 <= 32'b01111011011010000001000100101010;
op2 <= 32'b00100101101100011001110000100010;
#4;
op1 <= 32'b01101000111000001111011001111011;
op2 <= 32'b00011010000010000010011010100111;
#4;
op1 <= 32'b00010111001101100000011101110111;
op2 <= 32'b01001111011010010110111000101010;
#4;
op1 <= 32'b00000101000000001010111101000101;
op2 <= 32'b00000100000011100100001111001011;
#4;
op1 <= 32'b00110010101101000010111110100100;
op2 <= 32'b01111001000100100111000111001000;
#4;
op1 <= 32'b00100000100100011100001111011000;
op2 <= 32'b00101101101110011101001100000001;
#4;
op1 <= 32'b01001110100000000010011110101000;
op2 <= 32'b01100010101001101101110111011000;
#4;
op1 <= 32'b01111011111010001011001100111001;
op2 <= 32'b01010111000000001101111001000110;
#4;
op1 <= 32'b00101001010100110100110111010000;
op2 <= 32'b01001011100101100010101001000100;
#4;
op1 <= 32'b00010111101100111100100011001001;
op2 <= 32'b00000000101100011000100000001010;
#4;
op1 <= 32'b01000101100010000000001110001111;
op2 <= 32'b01110101111011111010001101100101;
#4;
op1 <= 32'b01110011110110110100111101010010;
op2 <= 32'b01101011001001111010011001110010;
#4;
op1 <= 32'b00100001010000100101101010111010;
op2 <= 32'b01011111100010111101001100001111;
#4;
op1 <= 32'b01001111110000011000001111011011;
op2 <= 32'b00010101000011101011110100100010;
#4;
op1 <= 32'b01111101100101010001011011011000;
op2 <= 32'b00001001101111111101000100111111;
#4;
op1 <= 32'b00101011010010011010011110100011;
op2 <= 32'b01111110010011010100111110001000;
#4;
op1 <= 32'b01011000101001110100010010100101;
op2 <= 32'b00110010111110010001010100010010;
#4;
op1 <= 32'b00000110111100110000110100010001;
op2 <= 32'b00101000001110110000100111001001;
#4;
op1 <= 32'b01110101001111000010001011100111;
op2 <= 32'b00011101011000011010010001011010;
#4;
op1 <= 32'b01100011010110001000111001001110;
op2 <= 32'b01010010100111101001100010011101;
#4;
op1 <= 32'b01001111111110001111011110111001;
op2 <= 32'b01000110001001100010100101110111;
#4;
op1 <= 32'b00111110001111101100101011101000;
op2 <= 32'b01111011100111110100110000111101;
#4;
op1 <= 32'b00101100101000110111010111011011;
op2 <= 32'b00110000101010010010100100111000;
#4;
op1 <= 32'b01011010000010111011101000100111;
op2 <= 32'b01100101010000010111101110001101;
#4;
op1 <= 32'b00000111111111000011101011011000;
op2 <= 32'b00011010010010010111000111110000;
#4;
op1 <= 32'b01110101110001100100110110101001;
op2 <= 32'b01001111000101001100111110010001;
#4;
op1 <= 32'b01100100000000100101000101111011;
op2 <= 32'b01000100011110100001101111110001;
#4;
op1 <= 32'b01010001100110001111101100001000;
op2 <= 32'b00111000111010000011000110101010;
#4;
op1 <= 32'b01111111101001001001111100010011;
op2 <= 32'b01101101111010111111010001010010;
#4;
op1 <= 32'b00101100111101000001111100011110;
op2 <= 32'b00100010010011010011011011100100;
#4;
op1 <= 32'b00011011010001111001111110100001;
op2 <= 32'b01010111101000010111000101111111;
#4;
op1 <= 32'b00001001010001111010001101001101;
op2 <= 32'b01001100100000110100110010010011;
#4;
op1 <= 32'b00110110110100010101111011111010;
op2 <= 32'b01000000111110110001101110100100;
#4;
op1 <= 32'b00100101000010111011100100011111;
op2 <= 32'b00110110011000010011010000001000;
#4;
op1 <= 32'b01010011001011000001010100001100;
op2 <= 32'b01101011011101110100100101100000;
#4;
op1 <= 32'b00000000100011110100111100000000;
op2 <= 32'b01011111110010000000101101010000;
#4;
op1 <= 32'b01101110100110111001110011101110;
op2 <= 32'b00010100111100100001011011101000;
#4;
op1 <= 32'b01011100010010101000111000000000;
op2 <= 32'b01001001011011011010100100001010;
#4;
op1 <= 32'b00001010000101110101011010001101;
op2 <= 32'b01111110001111010010010111101000;
#4;
op1 <= 32'b00110111111100011111100100101010;
op2 <= 32'b00110011010001001011110101000110;
#4;
op1 <= 32'b01100101011110001101011100010011;
op2 <= 32'b00100111110000101111010111111011;
#4;
op1 <= 32'b01010011110011111000000111000111;
op2 <= 32'b01011101001101100110011100010101;
#4;
op1 <= 32'b01000001101111110011001010010011;
op2 <= 32'b00010010000110101101001000101000;
#4;
op1 <= 32'b00101111110110111010100110011000;
op2 <= 32'b00000111001001101000001010000010;
#4;
op1 <= 32'b00011101011110110110001011100000;
op2 <= 32'b01111011110001001000010100100011;
#4;
op1 <= 32'b01001011000011110110000010100111;
op2 <= 32'b01110000010101100100001100000000;
#4;
op1 <= 32'b00111000110101001110000010000001;
op2 <= 32'b01100100111101100000011110000110;
#4;
op1 <= 32'b01100110100010111110101010011011;
op2 <= 32'b00011001110010010100100110010101;
#4;
op1 <= 32'b01010101000100111110100000110100;
op2 <= 32'b00001111010110111111111000111111;
#4;
op1 <= 32'b01000010110110101111000011101101;
op2 <= 32'b01000100010011011111100010100000;
#4;
op1 <= 32'b00110000111001110000010100110111;
op2 <= 32'b01111001000001000011011100100100;
#4;
op1 <= 32'b01011110010101110111001111000111;
op2 <= 32'b01101101100001100000110010011011;
#4;
op1 <= 32'b01001100101100111101110011110010;
op2 <= 32'b00100010111101010000011111011111;
#4;
op1 <= 32'b01111001111000000100010000111001;
op2 <= 32'b00010111000101110011011100101110;
#4;
op1 <= 32'b00101000010011010111110011011110;
op2 <= 32'b00001100100011001000110000100110;
#4;
op1 <= 32'b01010110100101000000101011000011;
op2 <= 32'b01000001111000110011111011001001;
#4;
op1 <= 32'b00000100100001000010101100111111;
op2 <= 32'b00110110111011100001001000110110;
#4;
op1 <= 32'b00110001111100000010111110010100;
op2 <= 32'b00101011011010100101110110111101;
#4;
op1 <= 32'b00011111110110000110011010111010;
op2 <= 32'b00100000010011010000010111110000;
#4;
op1 <= 32'b01001101111100010010110101010000;
op2 <= 32'b00010101000110110010001101001010;
#4;
op1 <= 32'b00111011110001100000111000010010;
op2 <= 32'b01001010000010101001111000010111;
#4;
op1 <= 32'b00101001011011011110110011001110;
op2 <= 32'b00111110110010100100110010101111;
#4;
op1 <= 32'b01010111001111100111011000100101;
op2 <= 32'b00110011100011011000111010010110;
#4;
op1 <= 32'b00000101100000111001000101000101;
op2 <= 32'b00101000110001110000010110001101;
#4;
op1 <= 32'b01110011011000000000011011111111;
op2 <= 32'b00011101100111000111001011101111;
#4;
op1 <= 32'b01100001001100001110101111001001;
op2 <= 32'b01010010100001110111001110111010;
#4;
op1 <= 32'b01001110001100110001001010001001;
op2 <= 32'b01000110100110100100110101101010;
#4;
op1 <= 32'b00111100010011100111010110000101;
op2 <= 32'b01111011100110000001011000110010;
#4;
op1 <= 32'b01101010010001000010100101010010;
op2 <= 32'b00110000011010010111011001001101;
#4;
op1 <= 32'b00010111110101011001111110010000;
op2 <= 32'b01100100111101100100111000110010;
#4;
op1 <= 32'b00000110000001000111100111001101;
op2 <= 32'b00011010010101111111000111001011;
#4;
op1 <= 32'b01110100001111100001111101001111;
op2 <= 32'b00001111100001100011100111101011;
#4;
op1 <= 32'b00100001101110101111100000001101;
op2 <= 32'b00000100000011011110110111000001;
#4;
op1 <= 32'b00001111111010110111001000110100;
op2 <= 32'b00111001010011110101000111010011;
#4;
op1 <= 32'b01111101110010001100000010001000;
op2 <= 32'b00101110000100111111101101100100;
#4;
op1 <= 32'b01101011101100100111011001011111;
op2 <= 32'b00100010110101101111100110010000;
#4;
op1 <= 32'b00011001110010001011000001001100;
op2 <= 32'b01011000000001111111000101111101;
#4;
op1 <= 32'b00000111011110100100001001000101;
op2 <= 32'b00001100110001010100110011011001;
#4;
op1 <= 32'b00110101100011111100101001111101;
op2 <= 32'b00000001110000001100001101001101;
#4;
op1 <= 32'b01100011100000100000001001110101;
op2 <= 32'b01110110111100011110011000111100;
#4;
op1 <= 32'b01010001010011110000011001101111;
op2 <= 32'b00101011101101101111010000011010;
#4;
op1 <= 32'b00111110100000100010111001110111;
op2 <= 32'b01011111111000110100100111011101;
#4;
op1 <= 32'b00101100100001000100111111001100;
op2 <= 32'b01010100101111110011011010110111;
#4;
op1 <= 32'b01011010110101010010100011000000;
op2 <= 32'b00001010010001010010101001110000;
#4;
op1 <= 32'b00001000100011001011000010001101;
op2 <= 32'b01111110101010001100101000011010;
#4;
op1 <= 32'b01110101101101011111001010100011;
op2 <= 32'b01110011001100010101011011101101;
#4;
op1 <= 32'b00100100100110001011101011101001;
op2 <= 32'b00101001000101111011011011001101;
#4;
op1 <= 32'b01010010000001101010110010001111;
op2 <= 32'b01011101010011101110111101110011;
#4;
op1 <= 32'b00000000000111010101001010010000;
op2 <= 32'b00010010011000110110011010001010;
#4;
op1 <= 32'b01101110001111110111100011110011;
op2 <= 32'b00000111100100101011011011110000;
#4;
op1 <= 32'b01011011100111110111010011110111;
op2 <= 32'b01111011111100001101001101111011;
#4;
op1 <= 32'b01001001101101001100000101010001;
op2 <= 32'b01110001000011111101101110110110;
#4;
op1 <= 32'b01110111100111001000111001001111;
op2 <= 32'b01100101111000101010110011011110;
#4;
op1 <= 32'b00100100110010101110010000100110;
op2 <= 32'b01011001110011010101001001100111;
#4;
op1 <= 32'b00010011000111110010100001101100;
op2 <= 32'b00001111100101000101111001000001;
#4;
op1 <= 32'b00000001000110010110001101111101;
op2 <= 32'b00000100011010010110001101101011;
#4;
op1 <= 32'b00101110111101011111100000100010;
op2 <= 32'b01111001001000000111000000111000;
#4;
op1 <= 32'b01011100101110110101101001010001;
op2 <= 32'b01101101111110011100010011101000;
#4;
op1 <= 32'b00001010010111001010110011010001;
op2 <= 32'b01100010101110010000110011111110;
#4;
op1 <= 32'b00111000001101110110010010011001;
op2 <= 32'b01010111011100101001011101101101;
#4;
op1 <= 32'b01100110101100100010001100010011;
op2 <= 32'b01001100111001110111001100000111;
#4;
op1 <= 32'b01010100110010100000001111010100;
op2 <= 32'b00000010001000010000001011111001;
#4;
op1 <= 32'b01000010010100111010100010111000;
op2 <= 32'b01110110110011011101100111010011;
#4;
op1 <= 32'b00110000001111011010101000100110;
op2 <= 32'b00101011100011101010010011011011;
#4;
op1 <= 32'b00011101110110011111101100100000;
op2 <= 32'b01100000010100110011000100110111;
#4;
op1 <= 32'b00001100010000100001110110110011;
op2 <= 32'b01010101011110101110001100111000;
#4;
op1 <= 32'b01111001001011101111100111100000;
op2 <= 32'b01001001010010101011011101001111;
#4;
op1 <= 32'b00100111111000111110000011101100;
op2 <= 32'b01111111001111111010011011010011;
#4;
op1 <= 32'b00010101001111110010111001100100;
op2 <= 32'b01110011011101111011110010101010;
#4;
op1 <= 32'b01000100001110111101101100101001;
op2 <= 32'b00101001100001010011001101111011;
#4;
op1 <= 32'b01110000111101111010001110011110;
op2 <= 32'b00011101011000110010001100010001;
#4;
op1 <= 32'b00011111000110001001011011101011;
op2 <= 32'b00010010011110100100101111100111;
#4;
op1 <= 32'b00001100100101100010011011111001;
op2 <= 32'b00000110111001100010110001110100;
#4;
op1 <= 32'b00111010101000010110100000111110;
op2 <= 32'b01111011111110100101110011101111;
#4;
op1 <= 32'b01101000001100111110010010001010;
op2 <= 32'b01110000100001100101100011001100;
#4;
op1 <= 32'b01010110101000000010011000101010;
op2 <= 32'b00100101111000111000000010110101;
#4;
op1 <= 32'b01000100000011001100010000000000;
op2 <= 32'b00011010011101100101110101001101;
#4;
op1 <= 32'b01110010001011110110011001000111;
op2 <= 32'b00001111100110010000111111001011;
#4;
op1 <= 32'b00100000011100010010001111111111;
op2 <= 32'b01000100110111111111001010011000;
#4;
op1 <= 32'b01001101110101100110101000011101;
op2 <= 32'b01111001001111010111000100110101;
#4;
op1 <= 32'b01111100001100011000101100010010;
op2 <= 32'b01101110101010110001111101110001;
#4;
op1 <= 32'b01101001100010011111100001101110;
op2 <= 32'b01100010101101010010101110001011;
#4;
op1 <= 32'b01010111011001010100010110001111;
op2 <= 32'b00011000000101010010010011110011;
#4;
op1 <= 32'b01000101001000001100010010011110;
op2 <= 32'b01001100011000011110000110101010;
#4;
op1 <= 32'b01110011100011010110000000001101;
op2 <= 32'b01000001111110100111001101000101;
#4;
op1 <= 32'b00100001001011100110011011110010;
op2 <= 32'b01110110100001111101011010101010;
#4;
op1 <= 32'b00001111001101000111011100010000;
op2 <= 32'b01101011101010000101010000110100;
#4;
op1 <= 32'b01111100100100101110010111111100;
op2 <= 32'b00011111101010001000110101111100;
#4;
op1 <= 32'b01101011000101001100110010000011;
op2 <= 32'b01010101010011000011010111011101;
#4;
op1 <= 32'b01011000101001000000000000100110;
op2 <= 32'b01001001111110111110110100001111;
#4;
op1 <= 32'b01000110010100000100001011101010;
op2 <= 32'b01111110101100011111100011110110;
#4;
op1 <= 32'b00110100001010001111011111011101;
op2 <= 32'b00110011011111110101001010111110;
#4;
op1 <= 32'b00100010010101010111001101100110;
op2 <= 32'b00101000101000101100110010101010;
#4;
op1 <= 32'b01010000100011001100111011101111;
op2 <= 32'b00011101111110110101011100111001;
#4;
op1 <= 32'b00111110000010110001110100010100;
op2 <= 32'b00010010001111000000001011100001;
#4;
op1 <= 32'b00101011110000000011110001000011;
op2 <= 32'b00000111001110111011001100100001;
#4;
op1 <= 32'b01011001101000011011001100011000;
op2 <= 32'b00111011111101101010001100111011;
#4;
op1 <= 32'b00000111111110101110100011110001;
op2 <= 32'b00110001010001101011111011001001;
#4;
op1 <= 32'b00110101100000101111110010101111;
op2 <= 32'b00100101110110001101000010101001;
#4;
op1 <= 32'b00100011110010110111001100001011;
op2 <= 32'b01011011011111010110100001001000;
#4;
op1 <= 32'b01010001000111110111011111000101;
op2 <= 32'b01001111011110111100011100011111;
#4;
op1 <= 32'b01111111011110100110001001100110;
op2 <= 32'b01000100111111100101011010101000;
#4;
op1 <= 32'b01101101000111001111011001111100;
op2 <= 32'b00111001010110000001110110011001;
#4;
op1 <= 32'b01011010101101000100011000000111;
op2 <= 32'b00101110001011010100110011011111;
#4;
op1 <= 32'b01001000100010101101101110100000;
op2 <= 32'b00100010111110000101000111111111;
#4;
op1 <= 32'b00110110000110000011011000000111;
op2 <= 32'b00010111100000101111101000101111;
#4;
op1 <= 32'b00100100110001110001000101110011;
op2 <= 32'b01001101000000010111101111001010;
#4;
op1 <= 32'b01010010000011100111101010111011;
op2 <= 32'b01000001100110110010111101111001;
#4;
op1 <= 32'b00000000100110110111000000101110;
op2 <= 32'b00110111001001101001110110100001;
#4;
op1 <= 32'b00101110001011000101000010100001;
op2 <= 32'b01101011100001010001101101011110;
#4;
op1 <= 32'b01011100100010110000111010001111;
op2 <= 32'b01100000111011110100111011010000;
#4;
op1 <= 32'b01001001110100010000111010100011;
op2 <= 32'b00010101001110111101100000001010;
#4;
op1 <= 32'b01110111110001010000000100100110;
op2 <= 32'b01001010001010000011100101110101;
#4;
op1 <= 32'b01100101100110111101110000100001;
op2 <= 32'b01111110110100110101100011010011;
#4;
op1 <= 32'b00010011001100100100010000010110;
op2 <= 32'b00110011100011011001110110000110;
#4;
op1 <= 32'b00000001011011100101010000110000;
op2 <= 32'b01101000101101111101100010000101;
#4;
op1 <= 32'b01101111100100111010100101000111;
op2 <= 32'b01011110000001111111001100111010;
#4;
op1 <= 32'b00011100101011110011011110011010;
op2 <= 32'b01010010000001001011000101010010;
#4;
op1 <= 32'b00001010100100100101010111110011;
op2 <= 32'b01000110111100110101110011100111;
#4;
op1 <= 32'b00111000110001001001011010110011;
op2 <= 32'b01111100000010000111001111110000;
#4;
op1 <= 32'b01100110100001011111001010111011;
op2 <= 32'b01110000111101101010101001101001;
#4;
op1 <= 32'b01010100100000001100101011010100;
op2 <= 32'b00100101110000111111011100011100;
#4;
op1 <= 32'b00000011001000111011010100110010;
op2 <= 32'b00011011011101101001001100011011;
#4;
op1 <= 32'b00110000000100010101111000001111;
op2 <= 32'b00001111101010100010110000010010;
#4;
op1 <= 32'b00011110011000001001001010100110;
op2 <= 32'b00000100110100001101011111001001;
#4;
op1 <= 32'b00001100100011101101011010000000;
op2 <= 32'b01111001110111111100101100000101;
#4;
op1 <= 32'b00111001101111101000000000101101;
op2 <= 32'b01101110001000100010000101010000;
#4;
op1 <= 32'b00100111111100000001011101110100;
op2 <= 32'b01100011100011100000010101000111;
#4;
op1 <= 32'b00010101100110100011010110010010;
op2 <= 32'b00011000000100011010000011111101;
#4;
op1 <= 32'b00000011100111011001011101011010;
op2 <= 32'b01001101000000101111110111011001;
#4;
op1 <= 32'b01110001101011011011111101010011;
op2 <= 32'b01000010001100011101111000001010;
#4;
op1 <= 32'b00011111000111101110010101010100;
op2 <= 32'b00110110100110111010110011100001;
#4;
op1 <= 32'b00001101000011100111111000111110;
op2 <= 32'b01101011100111110111000100110011;
#4;
op1 <= 32'b00111011001000000001100010011001;
op2 <= 32'b00100000100011001010110100100110;
#4;
op1 <= 32'b01101000110100010110101001001110;
op2 <= 32'b01010101000110001111001001001101;
#4;
op1 <= 32'b01010110011000000010000100100100;
op2 <= 32'b00001001111010101101101101100110;
#4;
op1 <= 32'b00000100000110101001100001011010;
op2 <= 32'b01111110100000110011100010011001;
#4;
op1 <= 32'b00110010011101100001001111010101;
op2 <= 32'b01110100000100000001101000000010;
#4;
op1 <= 32'b00100000010010000110000010100001;
op2 <= 32'b01101000101001010010011000111100;
#4;
op1 <= 32'b01001110011001011101100010111111;
op2 <= 32'b00011101110011011001100100100110;
#4;
op1 <= 32'b01111011111110101110001101001011;
op2 <= 32'b01010010011101001001100111110000;
#4;
op1 <= 32'b01101001110000101110010100010111;
op2 <= 32'b00000111000011011000000100001001;
#4;
op1 <= 32'b01011000011100000011001010010110;
op2 <= 32'b01111100110100101010010111100101;
#4;
op1 <= 32'b01000101111011111010000110010010;
op2 <= 32'b01110001001100000110011000010101;
#4;
op1 <= 32'b01110011110010100010011100011001;
op2 <= 32'b01100110000101111111100011100111;
#4;
op1 <= 32'b00100001111010000111110001001001;
op2 <= 32'b01011011011110110011100101000100;
#4;
op1 <= 32'b00001111111001011001110100001010;
op2 <= 32'b00010000011001100101110101101000;
#4;
op1 <= 32'b01111101100100101011010100100001;
op2 <= 32'b01000100110000110011101100011010;
#4;
op1 <= 32'b01101011001101100110001000101010;
op2 <= 32'b01111001100101001110111111110101;
#4;
op1 <= 32'b01011000111100111000000010111011;
op2 <= 32'b01101110011100001001000101111010;
#4;
op1 <= 32'b01000111000110100111011001100111;
op2 <= 32'b00100011011101101110101100011100;
#4;
op1 <= 32'b01110100110101111011011000010010;
op2 <= 32'b01011000000000101100111001011100;
#4;
op1 <= 32'b00100010100000010000011000111100;
op2 <= 32'b01001100111010000010111111101100;
#4;
op1 <= 32'b01010000010111110001110111001100;
op2 <= 32'b01000001101111000011101001110101;
#4;
op1 <= 32'b01111110100100101001101111011011;
op2 <= 32'b01110110111110101010010101001010;
#4;
op1 <= 32'b00101100010000110111111111001100;
op2 <= 32'b00101011111100110110000111111010;
#4;
op1 <= 32'b00011010010100011101110010011110;
op2 <= 32'b01100000101101110111000101110111;
#4;
op1 <= 32'b00000111100111001000001001101110;
op2 <= 32'b01010101001001000110101010001101;
#4;
op1 <= 32'b01110101111001110100100001110000;
op2 <= 32'b01001010011000000111111101110101;
#4;
op1 <= 32'b01100011100101101011011000010110;
op2 <= 32'b01111110111010010000100010111111;
#4;
op1 <= 32'b01010001001111010011001001111000;
op2 <= 32'b00110011110001001001001100111110;
#4;
op1 <= 32'b01111111111111110101110000001100;
op2 <= 32'b00101001100100000000101001111100;
#4;
op1 <= 32'b01101101011000001001001110001101;
op2 <= 32'b01011101101011010010000000001011;
#4;
op1 <= 32'b00011100000111110011100100000001;
op2 <= 32'b01010011101010111011011110110101;
#4;
op1 <= 32'b01001000110001101011100000010011;
op2 <= 32'b00000111010101001100010000100101;
#4;
op1 <= 32'b00110111001110110000111000011011;
op2 <= 32'b01111100100011110101010000100110;
#4;
op1 <= 32'b01100101000000101100101000011100;
op2 <= 32'b00110001010001100000101111100011;
#4;
op1 <= 32'b01010011001100001100101110001010;
op2 <= 32'b01100110100110101001110101000001;
#4;
op1 <= 32'b00000000011100000000011110011110;
op2 <= 32'b00011011000000011001100111100010;
#4;
op1 <= 32'b01101110110101100110101011001001;
op2 <= 32'b01010000010111100011001101000001;
#4;
op1 <= 32'b01011100010010101110000001010110;
op2 <= 32'b00000100101110110101001100100011;
#4;
op1 <= 32'b00001010110011110101001001101110;
op2 <= 32'b00111010010101011000100110000010;
#4;
op1 <= 32'b01110111110000101010110011010010;
op2 <= 32'b01101110010001000000011100001000;
#4;
op1 <= 32'b00100101111001110110001100101111;
op2 <= 32'b00100011011000011100111110111000;
#4;
op1 <= 32'b01010100000111000100100001111001;
op2 <= 32'b00011000100101011111011011011011;
#4;
op1 <= 32'b00000001111100110101110111110010;
op2 <= 32'b01001101001101010011011011011011;
#4;
op1 <= 32'b01101111100110001010101011000001;
op2 <= 32'b01000010010000001110010110001111;
#4;
op1 <= 32'b01011101000111101101110001110011;
op2 <= 32'b00110110100110101010001000101001;
#4;
op1 <= 32'b00001011001110110100001001110000;
op2 <= 32'b00101011101101000101001101101000;
#4;
op1 <= 32'b01111001010011111110101011001110;
op2 <= 32'b00100000101000101001101111100110;
#4;
op1 <= 32'b00100111001111011010010100011001;
op2 <= 32'b00010101110010100001111111000111;
#4;
op1 <= 32'b01010100010110010101111011100100;
op2 <= 32'b00001001100101010101010001000010;
#4;
op1 <= 32'b00000010011111110101100111101011;
op2 <= 32'b00111110111100100110000000001101;
#4;
op1 <= 32'b01110000111010001101110100101101;
op2 <= 32'b01110100010111001000000111110010;
#4;
op1 <= 32'b00011111010001000010110111001000;
op2 <= 32'b00101001110010011010111011100101;
#4;
op1 <= 32'b00001100101000011110010000100001;
op2 <= 32'b00011110010001110000111101101000;
#4;
op1 <= 32'b00111010010010100011100101100110;
op2 <= 32'b00010010111001010110100101101011;
#4;
op1 <= 32'b00101000011011010100011101001000;
op2 <= 32'b00000111110111000010011101010000;
#4;
op1 <= 32'b00010110001011111110000001011101;
op2 <= 32'b01111100100001001001100100110110;
#4;
op1 <= 32'b00000100000001111101110111100100;
op2 <= 32'b01110001101100111001000010111110;
#4;
op1 <= 32'b01110001101000111000011010101111;
op2 <= 32'b00100101111100100011101100011000;
#4;
op1 <= 32'b00011111101010100011011010110001;
op2 <= 32'b00011011010001010011111100001100;
#4;
op1 <= 32'b01001110010000110111010100101101;
op2 <= 32'b01010000101011000010101000000001;
#4;
op1 <= 32'b01111011110001010010110000101010;
op2 <= 32'b00000101010010111001000000001111;
#4;
op1 <= 32'b01101000111110001001101110100110;
op2 <= 32'b01111001010001000111011101000000;
#4;
op1 <= 32'b01010111010000011010011000111011;
op2 <= 32'b00101110110111110101001111101000;
#4;
op1 <= 32'b01000100110001110010001001101111;
op2 <= 32'b00100011000011111110100000000111;
#4;
op1 <= 32'b00110011010011111001001000101111;
op2 <= 32'b00011000101100101100100001010001;
#4;
op1 <= 32'b00100001000110100100110000001100;
op2 <= 32'b01001101101111000101101110011101;
#4;
op1 <= 32'b00001110110011010011001001111001;
op2 <= 32'b01000010001100010111100000000001;
#4;
op1 <= 32'b01111100110101101001011100010111;
op2 <= 32'b00110111010001011010000100010101;
#4;
op1 <= 32'b00101001101101101110111100111000;
op2 <= 32'b00101011011000000011100011101100;
#4;
op1 <= 32'b01011000100110001110001011101001;
op2 <= 32'b00100001000110001110000101010000;
#4;
op1 <= 32'b01000110000011000100001100111110;
op2 <= 32'b01010101011001000100010110100111;
#4;
op1 <= 32'b01110011111110101011100001110011;
op2 <= 32'b01001010011001110101011000000100;
#4;
op1 <= 32'b01100001111001001011000001101000;
op2 <= 32'b00111111011011111111011101101011;
#4;
op1 <= 32'b00010000010101000100001101110111;
op2 <= 32'b00110100101111111000110010100011;
#4;
op1 <= 32'b01111101100001101110001110100010;
op2 <= 32'b01101001000000110101110011001010;
#4;
op1 <= 32'b00101100000100011111111001000111;
op2 <= 32'b00011110101000110101101111011100;
#4;
op1 <= 32'b01011001000111110010010110110001;
op2 <= 32'b01010010101001110111111100011110;
#4;
op1 <= 32'b00000110111101111001110101000000;
op2 <= 32'b01000111100101110111001111100100;
#4;
op1 <= 32'b00110101001000100110001000100010;
op2 <= 32'b01111100011110011110111000101111;
#4;
op1 <= 32'b00100010110100110111011111100110;
op2 <= 32'b01110001000010101110100000110001;
#4;
op1 <= 32'b01010000100111010111011101001001;
op2 <= 32'b01100110011001110010101001000100;
#4;
op1 <= 32'b00111110011100010000011110110010;
op2 <= 32'b00011011000100111100111110011110;
#4;
op1 <= 32'b01101101000111101111110010100100;
op2 <= 32'b01010000101100011100101010100111;
#4;
op1 <= 32'b01011010110000100001100100000110;
op2 <= 32'b01000101001101101101110111100011;
#4;
op1 <= 32'b00001000100001100110011110011011;
op2 <= 32'b01111010000110011110111100011100;
#4;
op1 <= 32'b00110110001101101100001101000001;
op2 <= 32'b01101110101100010010101111001000;
#4;
op1 <= 32'b01100100010100011101001101110111;
op2 <= 32'b00100011110011010111100000010011;
#4;
op1 <= 32'b00010001110111001000101001101101;
op2 <= 32'b01011000001100110110011001010101;
#4;
op1 <= 32'b00000000000110100110101000001011;
op2 <= 32'b01001101101010011100100101011111;
#4;
op1 <= 32'b00101101101110010100101110001111;
op2 <= 32'b00000010001111011000000111011010;
#4;
op1 <= 32'b00011011100100111011100101010110;
op2 <= 32'b01110111001010100000110100110111;
#4;
op1 <= 32'b00001001101000111110011110101111;
op2 <= 32'b01101100000000110011111000010010;
#4;
op1 <= 32'b01110110111010010011100011100101;
op2 <= 32'b01100000010100111010001111001010;
#4;
op1 <= 32'b00100100111001111110011011000000;
op2 <= 32'b01010101011010011111101010100010;
#4;
op1 <= 32'b00010011000000111101000010111101;
op2 <= 32'b01001010100011011000000100010100;
#4;
op1 <= 32'b00000000111110101111001011010011;
op2 <= 32'b00111111011110011101000100100011;
#4;
op1 <= 32'b00101111000111101110110110000100;
op2 <= 32'b01110100100011011010010001011101;
#4;
op1 <= 32'b01011100110010001111110111110100;
op2 <= 32'b00101001011111101000101000111001;
#4;
op1 <= 32'b01001010110011101100000001001111;
op2 <= 32'b00011110010001111010100101001111;
#4;
op1 <= 32'b01111000011010001010101101100000;
op2 <= 32'b00010011000011001000010000110010;
#4;
op1 <= 32'b01100110001100111110000100110111;
op2 <= 32'b00000111101001011111100010010100;
#4;
op1 <= 32'b01010011111110110110010111000000;
op2 <= 32'b00111100011111100001100101001011;
#4;
op1 <= 32'b01000001110010110111001010010111;
op2 <= 32'b00110001000111111000011000100101;
#4;
op1 <= 32'b00110000000000100101011110100100;
op2 <= 32'b00100110100111010001010101110100;
#4;
op1 <= 32'b01011110001100011110010110110110;
op2 <= 32'b00011011100101110101111101100111;
#4;
op1 <= 32'b00001011011110101000111111101110;
op2 <= 32'b00010000000110000100100000011000;
#4;
op1 <= 32'b01111001111110100011010100010101;
op2 <= 32'b01000101100001111010011001110101;
#4;
op1 <= 32'b01100111011111011111100001011011;
op2 <= 32'b00111001111000011000001110100001;
#4;
op1 <= 32'b01010100101100011010001100101100;
op2 <= 32'b00101110001011111000111011110001;
#4;
op1 <= 32'b01000010110110001010111111101111;
op2 <= 32'b01100011011110011111101100110111;
#4;
op1 <= 32'b00110000111000100000111111001001;
op2 <= 32'b00011000010001101011000000111010;
#4;
op1 <= 32'b01011111001000001100101010100110;
op2 <= 32'b01001101110001111101101001011111;
#4;
op1 <= 32'b01001101001010101011000101100101;
op2 <= 32'b01000010111001110010100000011001;
#4;
op1 <= 32'b01111010010100100110110011001010;
op2 <= 32'b00110110110110110110001110101011;
#4;
op1 <= 32'b01101000011110001111100111001000;
op2 <= 32'b01101100000001111010000111001011;
#4;
op1 <= 32'b01010110011110000111100011010101;
op2 <= 32'b01100000111101110100111111011111;
#4;
op1 <= 32'b01000100100100010010011011011011;
op2 <= 32'b01010110000011110010000111011000;
#4;
op1 <= 32'b01110010001110110001000010011101;
op2 <= 32'b00001010110000010111010001011100;
#4;
op1 <= 32'b00011111110000101000111110001110;
op2 <= 32'b01111111011111111111011110011110;
#4;
op1 <= 32'b00001110100111110011010000001110;
op2 <= 32'b00110101000111000010011011001011;
#4;
op1 <= 32'b01111100001010011011100101010010;
op2 <= 32'b01101001101101001110000000101011;
#4;
op1 <= 32'b01101001100111100100101000011110;
op2 <= 32'b01011110001111101110000111111111;
#4;
op1 <= 32'b01010111010111101100110001010010;
op2 <= 32'b01010011000011011001000011001001;
#4;
op1 <= 32'b01000101101000101100101111011001;
op2 <= 32'b00001000000011111011001101001101;
#4;
op1 <= 32'b01110011010000101000000010111001;
op2 <= 32'b01111100110101010110000010000011;
#4;
op1 <= 32'b00100000110000111000011111111110;
op2 <= 32'b00110001010001110010010001011010;
#4;
op1 <= 32'b00001110110000100100111111101010;
op2 <= 32'b01100110010111100010101001101010;
#4;
op1 <= 32'b00111100100011001011101110011000;
op2 <= 32'b01011011001111010100111101111101;
#4;
op1 <= 32'b00101011000000100111010011010110;
op2 <= 32'b01010000100000010001110110110010;
#4;
op1 <= 32'b00011000101100011101000111110001;
op2 <= 32'b01000101010111001111100000000110;
#4;
op1 <= 32'b00000110010001011100110100111011;
op2 <= 32'b00111001110110010000000100110000;
#4;
op1 <= 32'b00110100001001011011000111101111;
op2 <= 32'b00101110110001001100010001010011;
#4;
op1 <= 32'b00100010001110100010011001101111;
op2 <= 32'b01100011101000101001000011001011;
#4;
op1 <= 32'b00001111100100010100110010010001;
op2 <= 32'b00011000000100010101101000000010;
#4;
op1 <= 32'b00111101101111110000000101100000;
op2 <= 32'b00001101010001100110111100101001;
#4;
op1 <= 32'b00101011101111010011001110001110;
op2 <= 32'b00000010011000001110011001101101;
#4;
op1 <= 32'b00011010000011110110111101111100;
op2 <= 32'b01110111101001100110000001101111;
#4;
op1 <= 32'b01001000000000100001110010101010;
op2 <= 32'b01101100101000100000101101101101;
#4;
op1 <= 32'b00110101001100110100011110100111;
op2 <= 32'b01100000101100000101100001010110;
#4;
op1 <= 32'b00100011001111110111111010100000;
op2 <= 32'b01010101101110110100100111010101;
#4;
op1 <= 32'b01010001001000100101101111110111;
op2 <= 32'b01001010101011011101111011101111;
#4;
op1 <= 32'b01111111010000010011001111100000;
op2 <= 32'b01111111111011110100010111111001;
#4;
op1 <= 32'b00101101011111011110010001000101;
op2 <= 32'b00110101000111010111001111011001;
#4;
op1 <= 32'b01011011001011010111000110100111;
op2 <= 32'b01101001111010011111010101110000;
#4;
op1 <= 32'b00001000110011011110011100001000;
op2 <= 32'b00011110010011011000010111011111;
#4;
op1 <= 32'b00110111001000101111100111000001;
op2 <= 32'b01010011100100001101011000101101;
#4;
op1 <= 32'b00100100101000101101001101111000;
op2 <= 32'b00001000010000110111101111010111;
#4;
op1 <= 32'b01010010011100100001100011110110;
op2 <= 32'b00111100111111001001110000110111;
#4;
op1 <= 32'b01000000100101011000010010001110;
op2 <= 32'b01110010000001001001101010111001;
#4;
op1 <= 32'b00101110011111010011000110010111;
op2 <= 32'b01100111000011000110110000100001;
#4;
op1 <= 32'b00011100001111010100000001010110;
op2 <= 32'b00011100000100110000000111011000;
#4;
op1 <= 32'b00001001111010011111011001000010;
op2 <= 32'b01010000010011001000011100110111;
#4;
op1 <= 32'b01110111110001101101011110011111;
op2 <= 32'b01000101010110101001100011010101;
#4;
op1 <= 32'b00100101011100010101111101011001;
op2 <= 32'b01111010000010001011111101111100;
#4;
op1 <= 32'b01010010111101111000110000100000;
op2 <= 32'b00101110100000001100011011010011;
#4;
op1 <= 32'b01000001000101101110100100010000;
op2 <= 32'b01100011100111010010100010011011;
#4;
op1 <= 32'b00101110111111011010011011010100;
op2 <= 32'b01011000100001100000010010100111;
#4;
op1 <= 32'b00011101001011000011100100110111;
op2 <= 32'b01001101101010110101111010100111;
#4;
op1 <= 32'b01001011000110000111001100111001;
op2 <= 32'b00000010110110011001010101000010;
#4;
op1 <= 32'b00111001000001101000100101001000;
op2 <= 32'b01110111101110100110010101001000;
#4;
op1 <= 32'b00100111001011000001010010010000;
op2 <= 32'b00101100100011010101111111001100;
#4;
op1 <= 32'b01010100110110110111010110111100;
op2 <= 32'b00100001010101111010110100000000;
#4;
op1 <= 32'b00000010010001001000101100110001;
op2 <= 32'b01010101110000000001100010000011;
#4;
op1 <= 32'b00110000011100001010100010111110;
op2 <= 32'b01001010111101100001000010010000;
#4;
op1 <= 32'b01011110000110100010100100010111;
op2 <= 32'b00111111101000100110001001011110;
#4;
op1 <= 32'b00001100110001100110101010010110;
op2 <= 32'b01110101011000100100001110000001;
#4;
op1 <= 32'b01111001101100111000011101011111;
op2 <= 32'b01101001001110111000110101010110;
#4;
op1 <= 32'b01101000000110010011100110010111;
op2 <= 32'b00011110110010011101110101010110;
#4;
op1 <= 32'b01010101010010011110000010110110;
op2 <= 32'b01010010111110110101001001100100;
#4;
op1 <= 32'b00000011101101001111110100100000;
op2 <= 32'b00001000001000111100110011000000;
#4;
op1 <= 32'b01110001001000010111110011111111;
op2 <= 32'b01111100100111111110101000011110;
#4;
op1 <= 32'b00011111010110100110100001011000;
op2 <= 32'b00110010000001111101100110000100;
#4;
op1 <= 32'b01001101000011100101000110100110;
op2 <= 32'b00100110101111011100111100100010;
#4;
op1 <= 32'b01111010111000101110001100111111;
op2 <= 32'b00011011011100001110110110010001;
#4;
op1 <= 32'b00101000110011011010001101001000;
op2 <= 32'b01010000100010110011001010001000;
#4;
op1 <= 32'b01010110010100001011010011100101;
op2 <= 32'b00000100111011010011000101000100;
#4;
op1 <= 32'b01000100111000110100101100111011;
op2 <= 32'b00111010011001011100010000000000;
#4;
op1 <= 32'b01110010101001100011111010100010;
op2 <= 32'b01101111001010001011011001100011;
#4;
op1 <= 32'b00100000010101100101001110100110;
op2 <= 32'b00100011111111101000111111000100;
#4;
op1 <= 32'b01001110100101001000101011010110;
op2 <= 32'b01011001000101011011110111010001;
#4;
op1 <= 32'b01111100011101101101010100000011;
op2 <= 32'b01001110010101100001000110100011;
#4;
op1 <= 32'b01101010010101011000001011111011;
op2 <= 32'b01000010111011111110000010011011;
#4;
op1 <= 32'b00011000011000110000100100011010;
op2 <= 32'b00111000000101001000101100010001;
#4;
op1 <= 32'b01000101111001110100001100000111;
op2 <= 32'b01101100011101001110111100100110;
#4;
op1 <= 32'b01110100010001101001011011011111;
op2 <= 32'b01100001111111111100111000111110;
#4;
op1 <= 32'b00100001001111000100111110111101;
op2 <= 32'b00010101101011110010100010000000;
#4;
op1 <= 32'b01001110111010001010000001111001;
op2 <= 32'b00001010010111101110010100110010;
#4;
op1 <= 32'b00111101011101100111010101110100;
op2 <= 32'b00000000001010000101111101100111;
#4;
op1 <= 32'b00101011000010011111011110101000;
op2 <= 32'b00110100011100111001111100011111;
#4;
op1 <= 32'b00011001010000000011110100111111;
op2 <= 32'b01101001111111100101110000111110;
#4;
op1 <= 32'b01000110111110000001000011000000;
op2 <= 32'b00011110100000111000101101001111;
#4;
op1 <= 32'b00110100000111101000000101010100;
op2 <= 32'b01010010101100101011111000110010;
#4;
op1 <= 32'b00100010100100001100001001011100;
op2 <= 32'b00001000000010011000000111111011;
#4;
op1 <= 32'b01010000100100000111110011001110;
op2 <= 32'b00111101000111010101101101111111;
#4;
op1 <= 32'b00111110010001000001010101101110;
op2 <= 32'b01110001100001100111001001101111;
#4;
op1 <= 32'b01101100100000000110111000100101;
op2 <= 32'b01100111001111000001100100110001;
#4;
op1 <= 32'b01011010101001010010010010000011;
op2 <= 32'b01011100010011001010100001011111;
#4;
op1 <= 32'b01001000100100001110111001100010;
op2 <= 32'b00010001001111011001110111110101;
#4;
op1 <= 32'b01110110000111000111011001111001;
op2 <= 32'b01000101100100100101110111100011;
#4;
op1 <= 32'b00100011000010001101111111000011;
op2 <= 32'b00111001110100011101001111010011;
#4;
op1 <= 32'b01010001100111111111111000111100;
op2 <= 32'b00101111001000011110001110110011;
#4;
op1 <= 32'b01111111011111100101100111011111;
op2 <= 32'b00100100000010001100011001111101;
#4;
op1 <= 32'b01101110000000111000010100000101;
op2 <= 32'b01011001101111010110011000110111;
#4;
op1 <= 32'b01011011001100101110011011111001;
op2 <= 32'b00001101111011111110100000010011;
#4;
op1 <= 32'b01001001000111100011100111110110;
op2 <= 32'b00000010110110111000100011010101;
#4;
op1 <= 32'b01110110110000111001100001110010;
op2 <= 32'b01110111100010100011010001011001;
#4;
op1 <= 32'b00100101011111010011101110110010;
op2 <= 32'b00101101000110011100111100001011;
#4;
op1 <= 32'b00010010010011010101101010011110;
op2 <= 32'b00100000110101110110001110001001;
#4;
op1 <= 32'b01000000110001011100111110001001;
op2 <= 32'b01010110100010101110110001001000;
#4;
op1 <= 32'b00101110000011111001101111101101;
op2 <= 32'b00001010101001101001010110000101;
#4;
op1 <= 32'b01011100110010111101111111100101;
op2 <= 32'b01000000010101111111101101100110;
#4;
op1 <= 32'b00001010001011001110000110110010;
op2 <= 32'b00110100111111010000001100011100;
#4;
op1 <= 32'b01110111101111000100101111110100;
op2 <= 32'b01101001011001111000011010110111;
#4;
op1 <= 32'b01100110001101111111001010011010;
op2 <= 32'b01011110110101101100111101111000;
#4;
op1 <= 32'b01010011100010101000100010110000;
op2 <= 32'b01010011010000001001010000100011;
#4;
op1 <= 32'b00000001101000110001101001000101;
op2 <= 32'b00001000001011101100110011000101;
#4;
op1 <= 32'b01101111010011010010000110100101;
op2 <= 32'b01111100110101101011000011111001;
#4;
op1 <= 32'b01011101010100000010101010111000;
op2 <= 32'b01110001111001011111101010010110;
#4;
op1 <= 32'b01001011001100001001010110010100;
op2 <= 32'b01100110111010011100010111111110;
#4;
op1 <= 32'b01111001100000011100000000101100;
op2 <= 32'b01011100000110111011111011000100;
#4;
op1 <= 32'b00100110111011010001000001111000;
op2 <= 32'b01010000011110001011011010110111;
#4;
op1 <= 32'b01010101001101101010111011010011;
op2 <= 32'b00000101111011010001100101100110;
#4;
op1 <= 32'b00000010101010001000111001000000;
op2 <= 32'b01111010000110111001000101101010;
#4;
op1 <= 32'b01110000100000010100110011010001;
op2 <= 32'b01101111001100100001111101011101;
#4;
op1 <= 32'b00011110001000011010111101001001;
op2 <= 32'b01100011101100001011111010001111;
#4;
op1 <= 32'b01001100101010011100010101100010;
op2 <= 32'b00011001010110101100001000110100;
#4;
op1 <= 32'b01111010100000101110111110001000;
op2 <= 32'b00001110010100100111110111010001;
#4;
op1 <= 32'b00101000001101001010011010001010;
op2 <= 32'b01000010111000101101111110011001;
#4;
op1 <= 32'b00010110001011110000000101001011;
op2 <= 32'b00110111111011111010000001110100;
#4;
op1 <= 32'b00000100010100010111001000101111;
op2 <= 32'b00101100111001001000101101110001;
#4;
op1 <= 32'b00110001011111011100100101101100;
op2 <= 32'b00100001001011011111100111000111;
#4;
op1 <= 32'b00011111110010000000000101110011;
op2 <= 32'b01010110011101100101101111010110;
#4;
op1 <= 32'b00001101000100000111100000101000;
op2 <= 32'b01001010110000101110101001001101;
#4;
op1 <= 32'b00111011001101111001001000101101;
op2 <= 32'b01111111111001011100100010110000;
#4;
op1 <= 32'b01101001011101010011100011001000;
op2 <= 32'b01110101001000101011101100100111;
#4;
op1 <= 32'b00010111010011010010110110111111;
op2 <= 32'b01101001111000001000010110100101;
#4;
op1 <= 32'b00000101000000011001010011101011;
op2 <= 32'b01011110101110111100001110110101;
#4;
op1 <= 32'b00110010110001010001001111110000;
op2 <= 32'b01010011100001000110000111111011;
#4;
op1 <= 32'b00100000100101010101111110010101;
op2 <= 32'b01001000000100000100111101011000;
#4;
op1 <= 32'b01001110010100011011010110111011;
op2 <= 32'b01111100110110000110000010010010;
#4;
op1 <= 32'b01111100011011101001001110011100;
op2 <= 32'b00110010010000110111101011000101;
#4;
op1 <= 32'b00101010000010110110100100011110;
op2 <= 32'b01100110101101101110101010100000;
#4;
op1 <= 32'b01011000100111111000010010000010;
op2 <= 32'b01011100010011101110110000111111;
#4;
op1 <= 32'b00000110100001001111111010111001;
op2 <= 32'b00010001001101101010110111110010;
#4;
op1 <= 32'b00110100000010100011001000101101;
op2 <= 32'b00000101110001111001101011000000;
#4;
op1 <= 32'b01100001101101111011110101111100;
op2 <= 32'b01111010010111001111000011010101;
#4;
op1 <= 32'b00001111010111010011111111101011;
op2 <= 32'b01101110111101001000000001100011;
#4;
op1 <= 32'b01111101100010000101110111100111;
op2 <= 32'b01100011111111000000101010110001;
#4;
op1 <= 32'b00101011100110101010101101111010;
op2 <= 32'b01011001001101101001000110010101;
#4;
op1 <= 32'b00011001011100011101100000011000;
op2 <= 32'b01001110010010111101100111001110;
#4;
op1 <= 32'b00000110111001100111110001110100;
op2 <= 32'b00000010100100010110000010110111;
#4;
op1 <= 32'b01110101010000000101110001011100;
op2 <= 32'b01110111100111101010001011010101;
#4;
op1 <= 32'b00100010110100111111011011110001;
op2 <= 32'b00101100100011001011001010011101;
#4;
op1 <= 32'b00010000101100010001111110001100;
op2 <= 32'b00100001011001000100011100101110;
#4;
op1 <= 32'b01111110110010100010001100100001;
op2 <= 32'b00010110011010001000000100000011;
#4;
op1 <= 32'b01101100111000010011000001001001;
op2 <= 32'b01001011110010100001111010101011;
#4;
op1 <= 32'b01011010011110101100111011001000;
op2 <= 32'b01000000011000000101101100000011;
#4;
op1 <= 32'b01001000100101001111001101001011;
op2 <= 32'b01110101011100100001111011110010;
#4;
op1 <= 32'b01110101111011010010110000110000;
op2 <= 32'b00101001101010011100001100111001;
#4;
op1 <= 32'b01100100000010001101001101001000;
op2 <= 32'b01011110110110011110101100111111;
#4;
op1 <= 32'b01010001110000001101010010100011;
op2 <= 32'b00010011011000100010110011001111;
#4;
op1 <= 32'b00111111101001110110100100100010;
op2 <= 32'b01001000010011011101110110111101;
#4;
op1 <= 32'b01101101010111000110101110110001;
op2 <= 32'b00111101000011010001110101011010;
#4;
op1 <= 32'b00011011101000010001011111100100;
op2 <= 32'b00110010010000101101000111100011;
#4;
op1 <= 32'b00001001000100001110011001101110;
op2 <= 32'b01100111000001100001001100100101;
#4;
op1 <= 32'b00110111101010100110000111010001;
op2 <= 32'b00011100011110001001010100111100;
#4;
op1 <= 32'b00100101011100001100010100011101;
op2 <= 32'b01010001001010110001000001111010;
#4;
op1 <= 32'b01010011000011001101100101110011;
op2 <= 32'b00000101101100001101111100111110;
#4;
op1 <= 32'b00000000100100000011100101100010;
op2 <= 32'b01111010011110110010101011010010;
#4;
op1 <= 32'b00101110010101001000010111000100;
op2 <= 32'b00101111000010110101000000100011;
#4;
op1 <= 32'b00011101000110001110011100100010;
op2 <= 32'b00100100110000100110001111111110;
#4;
op1 <= 32'b01001010101010010101001110010011;
op2 <= 32'b00011001011010010101001010001011;
#4;
op1 <= 32'b01111000110101001011011010101010;
op2 <= 32'b00001110100000110000111011010111;
#4;
op1 <= 32'b01100110010011101001101110110011;
op2 <= 32'b00000011000000100110011011100100;
#4;
op1 <= 32'b00010100011000101011111010011001;
op2 <= 32'b00111000000111000101111100101101;
#4;
op1 <= 32'b00000010010111001011001100010011;
op2 <= 32'b01101100111001101111010000011100;
#4;
op1 <= 32'b00110000000000100110101100000010;
op2 <= 32'b01100001100011000000110101100110;
#4;
op1 <= 32'b00011101001111111111001110101001;
op2 <= 32'b01010101110111010110100010101110;
#4;
op1 <= 32'b00001011101001001111100011011000;
op2 <= 32'b01001011011011110110000011001000;
#4;
op1 <= 32'b00111010001001000111010100010101;
op2 <= 32'b01000000101100001010011000010100;
#4;
op1 <= 32'b01100111011110101001000001110110;
op2 <= 32'b00110101000011111100011110010100;
#4;
op1 <= 32'b01010101000110101111010101011110;
op2 <= 32'b01101001110101000101111010011100;
#4;
op1 <= 32'b01000010110110111100001011110110;
op2 <= 32'b01011110100100110001100110101001;
#4;
op1 <= 32'b01110001011000010011010110011010;
op2 <= 32'b01010100000111101011110011100100;
#4;
op1 <= 32'b00011110110111100110000110001110;
op2 <= 32'b01001000011111010010110100011101;
#4;
op1 <= 32'b01001100111001100101100010100110;
op2 <= 32'b00111101101001010010100110011001;
#4;
op1 <= 32'b00111010100110001000101000101110;
op2 <= 32'b00110010100000000111011101110000;
#4;
op1 <= 32'b01101000110111100000100100101010;
op2 <= 32'b01100111110111100110101001101100;
#4;
op1 <= 32'b00010110110001111100111000010100;
op2 <= 32'b01011100011010110010111000000111;
#4;
op1 <= 32'b00000100101011000111011001111111;
op2 <= 32'b01010001100011000011101100110001;
#4;
op1 <= 32'b00110010010010010010001100110111;
op2 <= 32'b01000110000010101010000001000101;
#4;
op1 <= 32'b01100000010110011101110101001111;
op2 <= 32'b00111011000001100010101101101001;
#4;
op1 <= 32'b01001110000010110010010011111110;
op2 <= 32'b01101111100110001101100110000010;
#4;
op1 <= 32'b00111011111100111010111101100000;
op2 <= 32'b00100100110011100111100010101111;
#4;
op1 <= 32'b01101001111101010100010101011010;
op2 <= 32'b00011001101011011101101010100010;
#4;
op1 <= 32'b01010111000110010111111011111100;
op2 <= 32'b01001101110101000010010000000010;
#4;
op1 <= 32'b00000101111010111010000101010000;
op2 <= 32'b01000011110010001000110110111011;
#4;
op1 <= 32'b01110010101110010110001000110100;
op2 <= 32'b00110111010011001101101001010011;
#4;
op1 <= 32'b00100001010010010101001101011101;
op2 <= 32'b01101100111000101001110010001100;
#4;
op1 <= 32'b01001110101110101000101001101100;
op2 <= 32'b01100001011011011101110111111101;
#4;
op1 <= 32'b01111100111001010110111001111000;
op2 <= 32'b00010110100001100100011000001000;
#4;
op1 <= 32'b01101010100010000010101011100101;
op2 <= 32'b00001011011000011011011011001010;
#4;
op1 <= 32'b00011001000001011100000111110100;
op2 <= 32'b00000000111010100000011110001101;
#4;
op1 <= 32'b00000110000001111000111111110011;
op2 <= 32'b00110100100110010100110110101100;
#4;
op1 <= 32'b01110100110101011000110110111101;
op2 <= 32'b01101010100010101100110010111000;
#4;
op1 <= 32'b00100001100000001111010000110001;
op2 <= 32'b01011110010110100111010111101000;
#4;
op1 <= 32'b00010000000101010110000101111111;
op2 <= 32'b00010011101011011001110001101110;
#4;
op1 <= 32'b00111110000111010011101101100101;
op2 <= 32'b00001000101010011000011100010100;
#4;
op1 <= 32'b01101011110011100111001010001001;
op2 <= 32'b01111101011001100000011000111000;
#4;
op1 <= 32'b00011001010010111001111111110001;
op2 <= 32'b00110010000111100110110001000110;
#4;
op1 <= 32'b00000111010111010000111111100110;
op2 <= 32'b00100111000010010111000000101000;
#4;
op1 <= 32'b01110101101110101100010010000000;
op2 <= 32'b01011100101000000111110111010111;
#4;
op1 <= 32'b01100011101001110110110110101111;
op2 <= 32'b01010001010101111011101101010110;
#4;
op1 <= 32'b01010001011110010000100100111010;
op2 <= 32'b00000110010000100101000111011000;
#4;
op1 <= 32'b01111110101100100110011010000011;
op2 <= 32'b00111010011100111000001111111010;
#4;
op1 <= 32'b00101101100010101011110101011111;
op2 <= 32'b01110000010010111001111000111000;
#4;
op1 <= 32'b00011010111001100111011110100100;
op2 <= 32'b01100100100110001011011011001010;
#4;
op1 <= 32'b01001001011010110101011110001100;
op2 <= 32'b01011010010101010100000011100101;
#4;
op1 <= 32'b00110110011111010000110110101001;
op2 <= 32'b00001110010100110101011100100011;
#4;
op1 <= 32'b00100100001111110101001010100110;
op2 <= 32'b00000010111110011011100101110011;
#4;
op1 <= 32'b00010010100011100000110100111000;
op2 <= 32'b00111000010010000001101000111101;
#4;
op1 <= 32'b01000000010111001110001111010000;
op2 <= 32'b00101101000010110101001100000010;
#4;
op1 <= 32'b00101101011011101101010100010001;
op2 <= 32'b01100001001000011101000010000100;
#4;
op1 <= 32'b00011011101011111110110010100010;
op2 <= 32'b00010110010110100100010111000111;
#4;
op1 <= 32'b01001001100111111101110100111001;
op2 <= 32'b00001011010000111111011010010101;
#4;
op1 <= 32'b00110111110000011011100001101100;
op2 <= 32'b00000000010111101101000011101011;
#4;
op1 <= 32'b00100101101100011110100100011110;
op2 <= 32'b01110101100100100100010110101010;
#4;
op1 <= 32'b00010011011100110110010100001001;
op2 <= 32'b01101010001011010010001001001101;
#4;
op1 <= 32'b00000001011111101011100001001011;
op2 <= 32'b01011111010010101110010000101010;
#4;
op1 <= 32'b01101111011001010111100101010101;
op2 <= 32'b01010011111000110010010101110011;
#4;
op1 <= 32'b00011101100001000110000111101001;
op2 <= 32'b00001001100000100111110011100011;
#4;
op1 <= 32'b00001011000111001001111111101110;
op2 <= 32'b01111101110110001001111001000011;
#4;
op1 <= 32'b01111000111111101101110111001101;
op2 <= 32'b00110010110001110001111010011011;
#4;
op1 <= 32'b01100111010100100111011000101001;
op2 <= 32'b00101000000101010110101001101010;
#4;


end

always @(posedge clk) begin
    #4;
res_eth <= 32'b01110111101000010011011001111101;
#4;
res_eth <= 32'b00011010110010110100001100010101;
#4;
res_eth <= 32'b00111100100110001100010101010101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000010111110000101011111110110;
#4;
res_eth <= 32'b01100101011110010100001111101001;
#4;
res_eth <= 32'b00000110110111101010111000100110;
#4;
res_eth <= 32'b00101001111000010100001000101110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110001000101101101100000010100;
#4;
res_eth <= 32'b01010001100101100111011010100001;
#4;
res_eth <= 32'b00110101001101111000110001001101;
#4;
res_eth <= 32'b00010110101101110111011101110110;
#4;
res_eth <= 32'b00111011011011010110000000001010;
#4;
res_eth <= 32'b00011100100010110100000011000011;
#4;
res_eth <= 32'b00111111100111000100001101100011;
#4;
res_eth <= 32'b00100011001101011000000110101011;
#4;
res_eth <= 32'b01000101101110011010100000011110;
#4;
res_eth <= 32'b00101000111000000011101100110000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101101100111101100011000111000;
#4;
res_eth <= 32'b01010000111111010101100010111001;
#4;
res_eth <= 32'b01110100001001111001101010010101;
#4;
res_eth <= 32'b00010101100101101100001011111011;
#4;
res_eth <= 32'b01111001100010000001101001100111;
#4;
res_eth <= 32'b01011011101111011101110100100100;
#4;
res_eth <= 32'b01111111001010010111001111010110;
#4;
res_eth <= 32'b01100000100101101110100010010101;
#4;
res_eth <= 32'b00000101000001100010001111100000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00001000000111110100010011100010;
#4;
res_eth <= 32'b01101100101011001110011100010011;
#4;
res_eth <= 32'b01001111000001010100111110001001;
#4;
res_eth <= 32'b00110010001101001110000001011000;
#4;
res_eth <= 32'b00010100100001100000011000000010;
#4;
res_eth <= 32'b00110110111010100000101110100010;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00111101110101110000111111101110;
#4;
res_eth <= 32'b00011110101101100100001011010110;
#4;
res_eth <= 32'b01000011000110010011010101100001;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01001000000111011011100010111000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01001100110000000001111100111111;
#4;
res_eth <= 32'b01101111101001101000000001111010;
#4;
res_eth <= 32'b01010010110001101010111110111001;
#4;
res_eth <= 32'b00110101101011101111000111000101;
#4;
res_eth <= 32'b00011000001001011101100111110000;
#4;
res_eth <= 32'b00111010111111101101111101000010;
#4;
res_eth <= 32'b01011101100011001111110101101000;
#4;
res_eth <= 32'b00000001101110110100100101100010;
#4;
res_eth <= 32'b00100010010101001010100010100110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101000101001110111010011111100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101110100001111000001010101100;
#4;
res_eth <= 32'b01010000101011000111011000001001;
#4;
res_eth <= 32'b00110011101100011100010100011101;
#4;
res_eth <= 32'b01010110010010110011010001100011;
#4;
res_eth <= 32'b00111001100000001010101011000101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111111001010101111110110101000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01000100101011001011010011001100;
#4;
res_eth <= 32'b00100110111001100110011010110111;
#4;
res_eth <= 32'b00001010101111110110110111110001;
#4;
res_eth <= 32'b01101100011010001000111010001100;
#4;
res_eth <= 32'b01001110001000010001010010010101;
#4;
res_eth <= 32'b00110010100100000101101110111000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000000000011000;
#4;
res_eth <= 32'b01011001110101001000000010011011;
#4;
res_eth <= 32'b00000000000000000100001000101000;
#4;
res_eth <= 32'b01011111011011100111010100100110;
#4;
res_eth <= 32'b01000010001110101011111010011011;
#4;
res_eth <= 32'b00100100000000101000011101101000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00101010110010001011010010111111;
#4;
res_eth <= 32'b01001101101111101110000011100000;
#4;
res_eth <= 32'b01110000000000110110110100011010;
#4;
res_eth <= 32'b01010010101110010010010011000111;
#4;
res_eth <= 32'b00110110100010110010110011000000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00111011011110111001011101000111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000000000101100110110100011010;
#4;
res_eth <= 32'b00100100101101100011101001011110;
#4;
res_eth <= 32'b00000110010011101010001011000101;
#4;
res_eth <= 32'b00101000000100110111111011000011;
#4;
res_eth <= 32'b01001011010111000100111101111000;
#4;
res_eth <= 32'b00101110000011010101101001001010;
#4;
res_eth <= 32'b01010000110000111100001001110100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00010110011001011010110001001010;
#4;
res_eth <= 32'b00111001100010010100100110101010;
#4;
res_eth <= 32'b01011100000010101010010111101001;
#4;
res_eth <= 32'b00111110101100100000101001010001;
#4;
res_eth <= 32'b01100001010001000000000011110101;
#4;
res_eth <= 32'b01000100001001010111111111000001;
#4;
res_eth <= 32'b01100110100001010001011100101000;
#4;
res_eth <= 32'b01001001110001100111101010100010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110010111010111011101111000101;
#4;
res_eth <= 32'b01010100001001001100000010010011;
#4;
res_eth <= 32'b01111000001010010000101111011001;
#4;
res_eth <= 32'b01011010000101001110001000011011;
#4;
res_eth <= 32'b01111100101011000000111101100100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000011001111000001000111101010;
#4;
res_eth <= 32'b00100101011001010110010111101010;
#4;
res_eth <= 32'b01111111111110110000100101000010;
#4;
res_eth <= 32'b01101010101111011110110000101000;
#4;
res_eth <= 32'b00001101101010101101111011011100;
#4;
res_eth <= 32'b00110000001011010010101011110100;
#4;
res_eth <= 32'b01010011010010110101111000111110;
#4;
res_eth <= 32'b00110100111100110011111001000100;
#4;
res_eth <= 32'b01011000000010101110011111001110;
#4;
res_eth <= 32'b00111011000010000010001101001101;
#4;
res_eth <= 32'b01011101100001100000101100011011;
#4;
res_eth <= 32'b01000000011110001110101101100101;
#4;
res_eth <= 32'b00100011000111110001001011000000;
#4;
res_eth <= 32'b00000101110111011101100010010111;
#4;
res_eth <= 32'b01101001101011111110010100101011;
#4;
res_eth <= 32'b01001011100110000000000110010111;
#4;
res_eth <= 32'b00101110110110000110111000000010;
#4;
res_eth <= 32'b01010000011001011101001010001011;
#4;
res_eth <= 32'b00110100001100111001000010001010;
#4;
res_eth <= 32'b00010110001001111010011011111111;
#4;
res_eth <= 32'b00000000000000000000000010101000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111111000010101110010011101010;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01000100100100101101100100111111;
#4;
res_eth <= 32'b01111111110110111001101110011110;
#4;
res_eth <= 32'b01001000111000011100001000010001;
#4;
res_eth <= 32'b00101100101011110001000111100001;
#4;
res_eth <= 32'b01001111001100010111101000011011;
#4;
res_eth <= 32'b01110011000011110100011110111100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111000100011110100111110110101;
#4;
res_eth <= 32'b00011001101111000000111101010100;
#4;
res_eth <= 32'b00000000000000001000100100000101;
#4;
res_eth <= 32'b00100000100001110110001010001011;
#4;
res_eth <= 32'b01000011000011101011110110001100;
#4;
res_eth <= 32'b00100100010011001101101100101101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101010100000111000110111010111;
#4;
res_eth <= 32'b00001101010010001010011000100001;
#4;
res_eth <= 32'b00101111010101100110001010100111;
#4;
res_eth <= 32'b01010011011111011001011000001110;
#4;
res_eth <= 32'b01110101101010000011100001001100;
#4;
res_eth <= 32'b01011000100110100000011001110101;
#4;
res_eth <= 32'b01111011000001101111001101100001;
#4;
res_eth <= 32'b00011101100111011001001010111101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00100011010110110100101000111111;
#4;
res_eth <= 32'b01111111110100110011011010001110;
#4;
res_eth <= 32'b01101000010101000000011111010011;
#4;
res_eth <= 32'b01001100101001100101110111111111;
#4;
res_eth <= 32'b00101110000111010011100100100010;
#4;
res_eth <= 32'b01010000101111010101100011011110;
#4;
res_eth <= 32'b00110011111001000000000010100111;
#4;
res_eth <= 32'b00010101100110111111111100010001;
#4;
res_eth <= 32'b00000000000000000000100010111101;
#4;
res_eth <= 32'b01011011111111100101110010000000;
#4;
res_eth <= 32'b00111101101111001101010000100110;
#4;
res_eth <= 32'b00100001110010001011011011111001;
#4;
res_eth <= 32'b00000101001101010010100000110010;
#4;
res_eth <= 32'b00100111100111000110000100100100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101100110010011111110110011100;
#4;
res_eth <= 32'b01010000001111100010111101101100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010101011100110010100110110010;
#4;
res_eth <= 32'b00111000010000101111000001110101;
#4;
res_eth <= 32'b01011010010011100101010101011100;
#4;
res_eth <= 32'b00111101101101010001000011100100;
#4;
res_eth <= 32'b00011111100011001000000001011100;
#4;
res_eth <= 32'b01000010001101000100011000100110;
#4;
res_eth <= 32'b00100100110101000001101000100000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101001101110100110100010101001;
#4;
res_eth <= 32'b01001101101010110101010011011100;
#4;
res_eth <= 32'b00110000011100110110111111110100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00110110010100111000101001000111;
#4;
res_eth <= 32'b01011000110011110101110110111000;
#4;
res_eth <= 32'b00111011111000100010111000101110;
#4;
res_eth <= 32'b00011110011110000111001000110000;
#4;
res_eth <= 32'b01000001100010111011001001000001;
#4;
res_eth <= 32'b00100010101111111000110101001110;
#4;
res_eth <= 32'b00000110111000011100000110001000;
#4;
res_eth <= 32'b01101010000000101011010110000000;
#4;
res_eth <= 32'b00001010111010111110010010000010;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010010010000010000100111111011;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010111011110110110111000101011;
#4;
res_eth <= 32'b01111001110101111100110110101011;
#4;
res_eth <= 32'b01011100000110010010010100010110;
#4;
res_eth <= 32'b01111111001100101011000001101001;
#4;
res_eth <= 32'b00100001010011110101111010001100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01100110110110101100100101011011;
#4;
res_eth <= 32'b00001010100011110001011000100000;
#4;
res_eth <= 32'b00101100010000101011010011100110;
#4;
res_eth <= 32'b01010000000001001011110111001000;
#4;
res_eth <= 32'b01110010011100110001011000110100;
#4;
res_eth <= 32'b01010110000010011100100000100101;
#4;
res_eth <= 32'b01110111100100011000011100111011;
#4;
res_eth <= 32'b01011011000000000101001011011001;
#4;
res_eth <= 32'b00111101010010111000100011110010;
#4;
res_eth <= 32'b01011111100010001000010101110111;
#4;
res_eth <= 32'b01000010111010000111010111111010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01001000000110011010110001110011;
#4;
res_eth <= 32'b00101011100100000000110101010000;
#4;
res_eth <= 32'b01001101010010100111110011100010;
#4;
res_eth <= 32'b00110000001011000000100001010111;
#4;
res_eth <= 32'b00010011010011111100100011011010;
#4;
res_eth <= 32'b01110101101010010101000001010100;
#4;
res_eth <= 32'b00010111111010011110111111011111;
#4;
res_eth <= 32'b00000000000000000001101100110001;
#4;
res_eth <= 32'b00011101110001011101110001001010;
#4;
res_eth <= 32'b01000001000110111100101100001010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101001011001100000000010100100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101111101100000000011010100110;
#4;
res_eth <= 32'b00010001010000101111100010010101;
#4;
res_eth <= 32'b01110101001010110110111111101001;
#4;
res_eth <= 32'b01010111111010100100000100100100;
#4;
res_eth <= 32'b00111010011010101011100111111011;
#4;
res_eth <= 32'b00011011111010011111001001001011;
#4;
res_eth <= 32'b01111111000100101000111011000111;
#4;
res_eth <= 32'b00100010010101000110100010101111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01100110100000010001000101010100;
#4;
res_eth <= 32'b01001010101011101001111000101101;
#4;
res_eth <= 32'b00101100011010101101001010000011;
#4;
res_eth <= 32'b00001111101010101001001011011001;
#4;
res_eth <= 32'b01110010000101000011111010010001;
#4;
res_eth <= 32'b01010100001100000001010100100111;
#4;
res_eth <= 32'b00111000001111000010100010101000;
#4;
res_eth <= 32'b00011011010111110001010000010110;
#4;
res_eth <= 32'b00111101000001010101011110111000;
#4;
res_eth <= 32'b00011110111100100011110010101011;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01100110101100111011000001010101;
#4;
res_eth <= 32'b01001000100101111001101111011010;
#4;
res_eth <= 32'b00101011010101010000111010100000;
#4;
res_eth <= 32'b01001110100011111011101101111110;
#4;
res_eth <= 32'b01110000100100010101110000001111;
#4;
res_eth <= 32'b01010011001110010011101101100100;
#4;
res_eth <= 32'b00110110010000010011110110111010;
#4;
res_eth <= 32'b01011000111101111110111011001111;
#4;
res_eth <= 32'b00000000000000000101011110011101;
#4;
res_eth <= 32'b00011100111000111100100010101100;
#4;
res_eth <= 32'b00000001000010000100010011110100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101001001011011000110111101110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101110000101011011001111011001;
#4;
res_eth <= 32'b00010010000011100000111000111101;
#4;
res_eth <= 32'b01110011011101000111001010101000;
#4;
res_eth <= 32'b00010110110011000110110010100111;
#4;
res_eth <= 32'b00111001100001110000101111011111;
#4;
res_eth <= 32'b00011100100001101000111011001110;
#4;
res_eth <= 32'b01000000001101110101000111110100;
#4;
res_eth <= 32'b00100000101110010011011001110000;
#4;
res_eth <= 32'b00000100011001110110000011101101;
#4;
res_eth <= 32'b01100111010110010010011001011100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101100100101111001011111101000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01110010001000101010110100111111;
#4;
res_eth <= 32'b00010110000111100011111111011110;
#4;
res_eth <= 32'b00110111000001101010011100110111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000000000000011111110101001100;
#4;
res_eth <= 32'b00100001010000000111010010001110;
#4;
res_eth <= 32'b01000011010011000101011010110100;
#4;
res_eth <= 32'b01100101001100100101100101000111;
#4;
res_eth <= 32'b00000111110010000100101100000001;
#4;
res_eth <= 32'b01101011010011111110111110011111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101111100110100001111110011001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110101101100011011110111110111;
#4;
res_eth <= 32'b01011010000111101111010101110101;
#4;
res_eth <= 32'b01111100000111011111110110100110;
#4;
res_eth <= 32'b00011111011001111011101101011001;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01100100100111001100010000100011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101001101010011100010000110011;
#4;
res_eth <= 32'b01001100000101010101000011000101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010001001100000111001101101111;
#4;
res_eth <= 32'b00110100100001001111111011100010;
#4;
res_eth <= 32'b00010110110100101111010111101001;
#4;
res_eth <= 32'b00111001000011000101110000111100;
#4;
res_eth <= 32'b00011101100000110110011100011000;
#4;
res_eth <= 32'b00111111101011001001010111000011;
#4;
res_eth <= 32'b00100010101101011000010110010111;
#4;
res_eth <= 32'b00000100111000011100100000110010;
#4;
res_eth <= 32'b00100111001110110011100110100010;
#4;
res_eth <= 32'b01001010101000100000111100000100;
#4;
res_eth <= 32'b00101101100001100000011011100100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00110011100100101010100000010001;
#4;
res_eth <= 32'b01010110001000111111011110011111;
#4;
res_eth <= 32'b00111000010111101111010111001000;
#4;
res_eth <= 32'b00011011000101111101011110001110;
#4;
res_eth <= 32'b00111101111100110000110000010011;
#4;
res_eth <= 32'b00100000000000010101011011010101;
#4;
res_eth <= 32'b01000011001100001010001100101010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01001001010000001000010111100100;
#4;
res_eth <= 32'b01101011010010001000110100011001;
#4;
res_eth <= 32'b00001111010101010111101011101111;
#4;
res_eth <= 32'b01110010001011110100110110111010;
#4;
res_eth <= 32'b01010011001001111011101101101110;
#4;
res_eth <= 32'b00110110100101001001000110010101;
#4;
res_eth <= 32'b01011001100000100111001110010000;
#4;
res_eth <= 32'b00000000000000000101011000101101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01000001001111000100000010010011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000110001001000111100000100110;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101110011111111011001101010000;
#4;
res_eth <= 32'b01010011000010111100100111111011;
#4;
res_eth <= 32'b00110100111010010110100001011111;
#4;
res_eth <= 32'b00010111100110110101111101100011;
#4;
res_eth <= 32'b00000000000000000001100110001100;
#4;
res_eth <= 32'b00011101100000101010100111111110;
#4;
res_eth <= 32'b00111111010010100010111001101000;
#4;
res_eth <= 32'b01100011010101101111001101011011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00100111100011110110111110011000;
#4;
res_eth <= 32'b01001010010011100001111100100101;
#4;
res_eth <= 32'b01101100101101010000100100110111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01010101101100110001111000010001;
#4;
res_eth <= 32'b00000000000000000000000000010000;
#4;
res_eth <= 32'b00011011011110100111100010100110;
#4;
res_eth <= 32'b00111110100111100111011000100101;
#4;
res_eth <= 32'b01011111111111000001000011000110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00100101101111011111110001100010;
#4;
res_eth <= 32'b00001001111000010011111001011110;
#4;
res_eth <= 32'b00101100000010001000000100000101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01110000110001111111011101010011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01110110100111100000011101011001;
#4;
res_eth <= 32'b00011001010110001100011110110001;
#4;
res_eth <= 32'b00000000000000000001100111011111;
#4;
res_eth <= 32'b00011110100011001111001011000000;
#4;
res_eth <= 32'b01000010000000111110101100011000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000110101101110101011011100100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01001101000010110101010111101100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01010010101110000111010100000011;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010111101010000000110111110100;
#4;
res_eth <= 32'b00111010000001010100001011101100;
#4;
res_eth <= 32'b00011100110110001000101100111010;
#4;
res_eth <= 32'b00000000000011111111100011000101;
#4;
res_eth <= 32'b01100011010110101101011000001000;
#4;
res_eth <= 32'b01000100010110101111110111011101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101101010010111010100110001110;
#4;
res_eth <= 32'b01010000001010011011011110111001;
#4;
res_eth <= 32'b00110100000010100111011001111100;
#4;
res_eth <= 32'b01010110000101010100101100110010;
#4;
res_eth <= 32'b00111000000001111111001100011100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111101010100111000001000101010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000011110100011100001101110011;
#4;
res_eth <= 32'b01100101101001110010000010100001;
#4;
res_eth <= 32'b00000111101111101110010110001010;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01001101100001101110101001000111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110101100110110000001000110111;
#4;
res_eth <= 32'b01011001100111011011001110010001;
#4;
res_eth <= 32'b00000000000000000110010001100011;
#4;
res_eth <= 32'b01011111101110100011110011000010;
#4;
res_eth <= 32'b01000010000111001111010110111101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101001101110100101101111000011;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01101111110011100100001010111001;
#4;
res_eth <= 32'b00010010010000111100001111000001;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00010111010001100111010010001001;
#4;
res_eth <= 32'b00000000000000000000010001011000;
#4;
res_eth <= 32'b00011100101101011000100001001010;
#4;
res_eth <= 32'b00111110111000100101000010110001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000101011011100111101110010000;
#4;
res_eth <= 32'b00101000100010010010000001011111;
#4;
res_eth <= 32'b00001010111111001111000110111110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01110010110000000000011111011011;
#4;
res_eth <= 32'b01010100101110001001111011010010;
#4;
res_eth <= 32'b00111001000000111011001101111100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00111101110110011011000100010111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000011011111000011100011001011;
#4;
res_eth <= 32'b00100110000110000010010011100011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101100001101000000111110011000;
#4;
res_eth <= 32'b01001110011100000101011111101110;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010100110010010011110001010100;
#4;
res_eth <= 32'b00000000000000000000000000000101;
#4;
res_eth <= 32'b00011001000110011010100000111111;
#4;
res_eth <= 32'b00111100111000010110000010100100;
#4;
res_eth <= 32'b01011111001001111011100111000110;
#4;
res_eth <= 32'b01000001111010100100110100111001;
#4;
res_eth <= 32'b00100100100010111001111000100101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101010100101001010001110000111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01010010001111000111100100110100;
#4;
res_eth <= 32'b01110110011110101110101101101110;
#4;
res_eth <= 32'b00011000000111000010101111010000;
#4;
res_eth <= 32'b00111010101000101001111010111111;
#4;
res_eth <= 32'b00011101011111011100000010010001;
#4;
res_eth <= 32'b01000000010001101101100011110011;
#4;
res_eth <= 32'b01100011100011101000010001111100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01100111110101110101000010011101;
#4;
res_eth <= 32'b01001011000110001011111111001000;
#4;
res_eth <= 32'b00101111010000011011101011111101;
#4;
res_eth <= 32'b01010000001100000010110010010101;
#4;
res_eth <= 32'b01110010000010001011000110001011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01110110111001111000000111100011;
#4;
res_eth <= 32'b00011011000011000111001111101000;
#4;
res_eth <= 32'b00111110001011100100100000110011;
#4;
res_eth <= 32'b00100001100111111111010001011010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00100110100000000000001101011010;
#4;
res_eth <= 32'b00001000110000100001100101110001;
#4;
res_eth <= 32'b01101100011111010100110000100010;
#4;
res_eth <= 32'b01001111001010101111000000001100;
#4;
res_eth <= 32'b00110010000111001100011111010011;
#4;
res_eth <= 32'b01010101000101010110010111111110;
#4;
res_eth <= 32'b00000000000000000000000000011000;
#4;
res_eth <= 32'b00011010001000110000100100001101;
#4;
res_eth <= 32'b01111111110110010101111110110011;
#4;
res_eth <= 32'b01011111010111101001001010000111;
#4;
res_eth <= 32'b00000001101001101010001111011110;
#4;
res_eth <= 32'b00100100110111110000101010110000;
#4;
res_eth <= 32'b01000110111010011111111110110100;
#4;
res_eth <= 32'b01101011000100101011000001010010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110000011011000011100100000111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110100011001001010100100000100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00111010001101110111011001101100;
#4;
res_eth <= 32'b01011101001111110100101100100101;
#4;
res_eth <= 32'b00111111011001111001000001010100;
#4;
res_eth <= 32'b00100010011110000010111111100011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00100111001010100111000011000100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101101111101010010100101011111;
#4;
res_eth <= 32'b01010000000101000111110001111101;
#4;
res_eth <= 32'b01110100001111101111111001101000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00111001100001111000101111010101;
#4;
res_eth <= 32'b01011100000010011111110101010000;
#4;
res_eth <= 32'b00000000000001110101000011000100;
#4;
res_eth <= 32'b01100001101000010000000101100111;
#4;
res_eth <= 32'b01000011011011110100100111010001;
#4;
res_eth <= 32'b00100111001001011111101100100000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01101100010011100010011010000011;
#4;
res_eth <= 32'b00001110110100111001110101011000;
#4;
res_eth <= 32'b01110001101001110001000110001011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110101011101111110010011110110;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111011111111101010010001000101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000001010101000100111011111110;
#4;
res_eth <= 32'b00100101010101111100110000110111;
#4;
res_eth <= 32'b01000111110111110110101111001111;
#4;
res_eth <= 32'b01101010001000011011100111100011;
#4;
res_eth <= 32'b01001100001000101011111110001001;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010011001001011101001101110110;
#4;
res_eth <= 32'b01110110100001100010100011101101;
#4;
res_eth <= 32'b01010110101000011001100011110101;
#4;
res_eth <= 32'b01111010011011010111000110110000;
#4;
res_eth <= 32'b00011101110110000000011000111110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101000111111101010001110010111;
#4;
res_eth <= 32'b01001011000010101100000100101101;
#4;
res_eth <= 32'b01111111111001001001111100010011;
#4;
res_eth <= 32'b00001111110000111011000101000011;
#4;
res_eth <= 32'b00110011011110111100011111001001;
#4;
res_eth <= 32'b00010110010011001100100010001111;
#4;
res_eth <= 32'b00111000010011010101111010111010;
#4;
res_eth <= 32'b00011011111101011101010000110100;
#4;
res_eth <= 32'b01111111001001100011100110100001;
#4;
res_eth <= 32'b00100000110111111111100000011010;
#4;
res_eth <= 32'b01000100000100110010100001000101;
#4;
res_eth <= 32'b01100110001111000000101100110110;
#4;
res_eth <= 32'b01001000110111111010001010011110;
#4;
res_eth <= 32'b00101011101110011111010110101011;
#4;
res_eth <= 32'b01001101101111011000001000010110;
#4;
res_eth <= 32'b01110001100100111101100111010010;
#4;
res_eth <= 32'b00010100011001110100001011000100;
#4;
res_eth <= 32'b00000000000000000000000000100100;
#4;
res_eth <= 32'b01011001110000001111101001110000;
#4;
res_eth <= 32'b01111011111100000000000010100100;
#4;
res_eth <= 32'b01011110010011001001010111111110;
#4;
res_eth <= 32'b01000000110111000000011011010110;
#4;
res_eth <= 32'b00100100111111100011010100010011;
#4;
res_eth <= 32'b01000111101100000010011110010000;
#4;
res_eth <= 32'b01101010011011101010000011100110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110000001011000010011111111011;
#4;
res_eth <= 32'b01010001100001000111100010010101;
#4;
res_eth <= 32'b00000000000000000000000000000010;
#4;
res_eth <= 32'b01011001000000110110100111011010;
#4;
res_eth <= 32'b00000000000000000011110101110101;
#4;
res_eth <= 32'b00011101110110111110001101110000;
#4;
res_eth <= 32'b00000000101011010100111101001000;
#4;
res_eth <= 32'b00100011100100100010011110101110;
#4;
res_eth <= 32'b01000110010101100111101111001000;
#4;
res_eth <= 32'b00101000101111000000010000011111;
#4;
res_eth <= 32'b01001011010100101010001001001111;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010001100010001110100011011000;
#4;
res_eth <= 32'b01110100001110110011100010100011;
#4;
res_eth <= 32'b01010101010101111101111010011010;
#4;
res_eth <= 32'b01111000011101010100111101011011;
#4;
res_eth <= 32'b01011011001100101110010001000010;
#4;
res_eth <= 32'b00111101010011011000100010010101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01000100010001110101111011001110;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00001001101111101010110010011001;
#4;
res_eth <= 32'b01101100011010000001011101100011;
#4;
res_eth <= 32'b01001111000101011101110011101101;
#4;
res_eth <= 32'b00110010010101010010010010010000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000000000110110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111101100100111111001111111010;
#4;
res_eth <= 32'b01011110111001110010100110000110;
#4;
res_eth <= 32'b01000001110001011010011110100001;
#4;
res_eth <= 32'b00100101101001000010101110110010;
#4;
res_eth <= 32'b01000111101110011000010111011100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00001110001101010000011010011101;
#4;
res_eth <= 32'b01101111110110011011100110100101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00110110010110110111011110011100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111011010010110010011000111100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111111001000101011101000000001;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01101000100110100010011011101000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101101100111111000010000010110;
#4;
res_eth <= 32'b01010000001011011100100110010011;
#4;
res_eth <= 32'b01110100001000010000110110110001;
#4;
res_eth <= 32'b00010111011111100001110110000010;
#4;
res_eth <= 32'b01111001101010100011001000110100;
#4;
res_eth <= 32'b00011100010100110101110100001001;
#4;
res_eth <= 32'b00111110101100111101001111100011;
#4;
res_eth <= 32'b00100010001111100011110101001100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01100111101010101001100101010000;
#4;
res_eth <= 32'b01001001001110010000001010101000;
#4;
res_eth <= 32'b00101110010000110111110101000110;
#4;
res_eth <= 32'b01001110110110111011100000000001;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01110111000111011101101001100101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111101000011100101001001011100;
#4;
res_eth <= 32'b00011111000001110111011110100110;
#4;
res_eth <= 32'b01000010010100011011110111100101;
#4;
res_eth <= 32'b00100101110100101111001011011110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110000000001011001001010010100;
#4;
res_eth <= 32'b01010010000011011101101010000110;
#4;
res_eth <= 32'b01110110000010100100111101110101;
#4;
res_eth <= 32'b01011000001110010001010100001111;
#4;
res_eth <= 32'b00111011011011010101001011111100;
#4;
res_eth <= 32'b01011100110000010111000000111010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01100011001000010110010000000011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101000001010001000010110000010;
#4;
res_eth <= 32'b00001011100001111011110110101100;
#4;
res_eth <= 32'b00101111000010100011111011011110;
#4;
res_eth <= 32'b00010000110011000101010111010110;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010110000110111100100100110011;
#4;
res_eth <= 32'b00000000000000000000001100001011;
#4;
res_eth <= 32'b00011011110111011101111111101111;
#4;
res_eth <= 32'b00111111110010010110001110010010;
#4;
res_eth <= 32'b01100001000111001101011001111000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01100111000001001000001000011110;
#4;
res_eth <= 32'b01001001011101000001001011101001;
#4;
res_eth <= 32'b00101100000001101011000100111101;
#4;
res_eth <= 32'b00001110000110111100000001100001;
#4;
res_eth <= 32'b00110010010010010110000000011011;
#4;
res_eth <= 32'b01010100001011001011110101110110;
#4;
res_eth <= 32'b00000000000000000000000001100101;
#4;
res_eth <= 32'b01011010001100110011000010011111;
#4;
res_eth <= 32'b01111110000000011111110101100111;
#4;
res_eth <= 32'b00011111100110010110011000011110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000111010001010011101001100010;
#4;
res_eth <= 32'b00101010101010110010011111000001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101111001101011010010000010010;
#4;
res_eth <= 32'b00010010000010110001110010110001;
#4;
res_eth <= 32'b01110101010100011001001000101110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111010110001010010110110100011;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00000000011000001010000101111100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01000110111110011011110001000001;
#4;
res_eth <= 32'b01101000011100010100101111001101;
#4;
res_eth <= 32'b01001100000001010011000111110101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00010001001000010100011001000000;
#4;
res_eth <= 32'b01110100011100010110111111110110;
#4;
res_eth <= 32'b00010110010000010100000001001111;
#4;
res_eth <= 32'b00111001001100010111111011010101;
#4;
res_eth <= 32'b00011100001011111111001101111000;
#4;
res_eth <= 32'b01111110011110100011101010101000;
#4;
res_eth <= 32'b00100000110011011001111001100001;
#4;
res_eth <= 32'b01000011000111100111110001001000;
#4;
res_eth <= 32'b01100111000010101000010000101000;
#4;
res_eth <= 32'b01001001100000010100010000110101;
#4;
res_eth <= 32'b00101100101110001001100000010010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110001010101110111010011010100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01110111101001010001111010100010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111101111001000010010111011101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101011000101001111101110100011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101111111010100000101110011011;
#4;
res_eth <= 32'b01010010101001000000110011010101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00011000101110011101110100100001;
#4;
res_eth <= 32'b00111011100101100110000110111001;
#4;
res_eth <= 32'b00011101010010010000100101100101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000101100100010100011101110110;
#4;
res_eth <= 32'b01111111111111110101110000001100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110000010101011001101010101100;
#4;
res_eth <= 32'b00010000101001010010100010110001;
#4;
res_eth <= 32'b01110100010100010111010010111011;
#4;
res_eth <= 32'b01010110110010100101110011001001;
#4;
res_eth <= 32'b01111010010101011000111000010101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00100001100101000111001111000001;
#4;
res_eth <= 32'b00000101101011001110111011110010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00001001110011000001100111101100;
#4;
res_eth <= 32'b00101101001101110001100111000100;
#4;
res_eth <= 32'b00001111101011000100010110010010;
#4;
res_eth <= 32'b01110010011001100001000111101110;
#4;
res_eth <= 32'b01010100001111111110101001111100;
#4;
res_eth <= 32'b00000000000000000000000000100001;
#4;
res_eth <= 32'b01011010100001000001000100110100;
#4;
res_eth <= 32'b00000000000000100101011011101111;
#4;
res_eth <= 32'b00011110011111011001011110001100;
#4;
res_eth <= 32'b00000001111100011100001011001111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00001001100110101000110111111001;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00001101101101010011100010011110;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010011001101100011000111100100;
#4;
res_eth <= 32'b00110110001111101001100111110000;
#4;
res_eth <= 32'b01011000000110101011101100010001;
#4;
res_eth <= 32'b00000000000000000010000011001010;
#4;
res_eth <= 32'b01011111100000110111001011001100;
#4;
res_eth <= 32'b01000001100111001100100011111010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000110101010001110111101000110;
#4;
res_eth <= 32'b00101000010111111110000101110001;
#4;
res_eth <= 32'b00001100100100001111011000010001;
#4;
res_eth <= 32'b00101111011000110000111000100001;
#4;
res_eth <= 32'b00010001100011100100000000010110;
#4;
res_eth <= 32'b01110100101001011010100101001011;
#4;
res_eth <= 32'b00010101101000000011100111111110;
#4;
res_eth <= 32'b00111010001101101001101010010011;
#4;
res_eth <= 32'b01011011111110100010010000011010;
#4;
res_eth <= 32'b01111110111000101001000010101110;
#4;
res_eth <= 32'b01100001110101100101110110110111;
#4;
res_eth <= 32'b00000101100111101101001011110010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00001011001110100101001010010100;
#4;
res_eth <= 32'b01101100010100000100000100111010;
#4;
res_eth <= 32'b00001111000100100111110111011001;
#4;
res_eth <= 32'b01110010000111101000100010001000;
#4;
res_eth <= 32'b01010100011001010111110011011110;
#4;
res_eth <= 32'b01110111100011100011000010100010;
#4;
res_eth <= 32'b00011010000010110010101011100101;
#4;
res_eth <= 32'b01111110010111001101010100010001;
#4;
res_eth <= 32'b01100000100010101010011000000110;
#4;
res_eth <= 32'b01000011001000011010001011101010;
#4;
res_eth <= 32'b01100101011111001111100010000011;
#4;
res_eth <= 32'b01001000101010000110100011000001;
#4;
res_eth <= 32'b00101010100110101000110011110011;
#4;
res_eth <= 32'b00001101100011000010011001000011;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010011010001000100000101100111;
#4;
res_eth <= 32'b00110110001010000000111010011000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111010110100111111010000001111;
#4;
res_eth <= 32'b00011110000100011011100011011101;
#4;
res_eth <= 32'b00000000111101001110001100110010;
#4;
res_eth <= 32'b01100100001011111101110110110111;
#4;
res_eth <= 32'b01000110110001111101100001111110;
#4;
res_eth <= 32'b00101001101000010100000000111010;
#4;
res_eth <= 32'b01001011111111110110101110111101;
#4;
res_eth <= 32'b00101110011010010011110110100101;
#4;
res_eth <= 32'b01010000111110011000011111001011;
#4;
res_eth <= 32'b00110011011111011000110110001110;
#4;
res_eth <= 32'b00010111000111111111010101011000;
#4;
res_eth <= 32'b00111010010100100110000110010100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01100001110111111011100111011110;
#4;
res_eth <= 32'b01000011011100111010001101110110;
#4;
res_eth <= 32'b01100110110100111001011111000011;
#4;
res_eth <= 32'b00001001101011110111001111010100;
#4;
res_eth <= 32'b01101101011110110000110101011111;
#4;
res_eth <= 32'b01010000100110100010000011001111;
#4;
res_eth <= 32'b01110001101101000101010011111101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01110111111100000000101000011011;
#4;
res_eth <= 32'b01011011001000100100111111001010;
#4;
res_eth <= 32'b00111101100011010101110010001101;
#4;
res_eth <= 32'b01011111110000101000100100101111;
#4;
res_eth <= 32'b00000100010000100011011110110001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101010111101100110100100010110;
#4;
res_eth <= 32'b00001110001101101100001111000111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00010010100110000001101001111010;
#4;
res_eth <= 32'b00110101101010001010000101111110;
#4;
res_eth <= 32'b01011000010100000010010001100100;
#4;
res_eth <= 32'b00111100000000111001100000000100;
#4;
res_eth <= 32'b00011110100110010111110010110011;
#4;
res_eth <= 32'b00000000101001111010101111100010;
#4;
res_eth <= 32'b00100011011111101011011010011010;
#4;
res_eth <= 32'b01000110011011000110101100110111;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00001011100101000000111000000000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010010001110100111000010100101;
#4;
res_eth <= 32'b01110101001001001011011111100100;
#4;
res_eth <= 32'b01010110011101101111111000111111;
#4;
res_eth <= 32'b00111001100011000001100010111001;
#4;
res_eth <= 32'b01011100010111001000101100010010;
#4;
res_eth <= 32'b01111111111011110100010111111001;
#4;
res_eth <= 32'b00100011000111000010011111100011;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01001011001110000110100110101100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01001111111011101110010001001101;
#4;
res_eth <= 32'b01110011000110101110010101101110;
#4;
res_eth <= 32'b01010110000010101110001000010000;
#4;
res_eth <= 32'b00000000000000000000000011011001;
#4;
res_eth <= 32'b00011010101110101110101111010000;
#4;
res_eth <= 32'b01111101101010011100101001010011;
#4;
res_eth <= 32'b01100000000000001110111100110010;
#4;
res_eth <= 32'b01000001111110010000110010100101;
#4;
res_eth <= 32'b01100101001110010100100110111101;
#4;
res_eth <= 32'b01001000000001001100100111101111;
#4;
res_eth <= 32'b00101011011001101001001111001010;
#4;
res_eth <= 32'b00001110100000011001001010001110;
#4;
res_eth <= 32'b01110001010000111110100111110001;
#4;
res_eth <= 32'b00010100001111100000111101110000;
#4;
res_eth <= 32'b00110110101110001110010000101111;
#4;
res_eth <= 32'b00011000100100110111101100110110;
#4;
res_eth <= 32'b00111011111001110101000110111000;
#4;
res_eth <= 32'b01011110010000111001001001111010;
#4;
res_eth <= 32'b01000010101011110101111001101010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000111011100011010010101100011;
#4;
res_eth <= 32'b01101000110001100011000001001011;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00010001111001111100110100110011;
#4;
res_eth <= 32'b00110100010100110000101011011101;
#4;
res_eth <= 32'b01010110110101011000011110011000;
#4;
res_eth <= 32'b00111001110111111010000001111110;
#4;
res_eth <= 32'b00011011110000010101111110100010;
#4;
res_eth <= 32'b00111111110011000000000001010001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000100110101010001111101011100;
#4;
res_eth <= 32'b01101000001011011100010111100101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101101110010000001000010011100;
#4;
res_eth <= 32'b00010001000000111011110010011000;
#4;
res_eth <= 32'b01110010110111010100001111101101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000000000100000;
#4;
res_eth <= 32'b00011001110010101000101101101110;
#4;
res_eth <= 32'b00000000000000100110110111100011;
#4;
res_eth <= 32'b00100000000000110100101111010110;
#4;
res_eth <= 32'b01000011101111110000001000001001;
#4;
res_eth <= 32'b00100101111111101110111100100000;
#4;
res_eth <= 32'b01000111010111010101011101011111;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01001110001100011010000001011101;
#4;
res_eth <= 32'b01110000010011011111010110111100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01110111100001000000010110110110;
#4;
res_eth <= 32'b00011010010101101011001011010111;
#4;
res_eth <= 32'b01111100001100101110100111100110;
#4;
res_eth <= 32'b00011101011000000101111111011111;
#4;
res_eth <= 32'b01000001010010100101101001100100;
#4;
res_eth <= 32'b01100100000001111110010011110100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00101001101001111010011111010001;
#4;
res_eth <= 32'b00001100100001111011000000101000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00010011000110000010010101111100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010111110101101011000011100110;
#4;
res_eth <= 32'b00000000000000000000000101110110;
#4;
res_eth <= 32'b01011101101011000000000100111111;
#4;
res_eth <= 32'b00000000001010101011011101001010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01100111010100000110110101011100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01110010101000010100000010110110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110111111001100101000100100111;
#4;
res_eth <= 32'b00011011101010010011000111111001;
#4;
res_eth <= 32'b00111101010011001101101110111110;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000010010111110100000110111001;
#4;
res_eth <= 32'b00100110100100010001001011100000;
#4;
res_eth <= 32'b01001001010101110101000110101111;
#4;
res_eth <= 32'b00101011101000000001100011001111;
#4;
res_eth <= 32'b00001110101000111100111111100101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00010011001011000111100010111100;
#4;
res_eth <= 32'b00110110110000000111100100100100;
#4;
res_eth <= 32'b00011000010110111111111010001111;
#4;
res_eth <= 32'b01111111111001011100100010110000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000001101100111111001100100100;
#4;
res_eth <= 32'b00100100001111100001010110101111;
#4;
res_eth <= 32'b01000110110010111101001101101011;
#4;
res_eth <= 32'b00101001001010000110100000011111;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01101111001101100010110011011010;
#4;
res_eth <= 32'b01010001010001110011100100000001;
#4;
res_eth <= 32'b01110101100000001110111111010110;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000011010111100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00111110110100110100111111100010;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000101010111001001101110111100;
#4;
res_eth <= 32'b00101000010000001001010000011110;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00001111111010001111110111011111;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01010101101101111001010110110100;
#4;
res_eth <= 32'b01111001001100011100101100010100;
#4;
res_eth <= 32'b01011011010110111100111000011001;
#4;
res_eth <= 32'b01111110100011001101111111111110;
#4;
res_eth <= 32'b01100000000111010100011100001001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00100101101010100101110101111000;
#4;
res_eth <= 32'b01001000100001101010000000110010;
#4;
res_eth <= 32'b01101010111100110000000100101100;
#4;
res_eth <= 32'b00001110011101010011000001011100;
#4;
res_eth <= 32'b00110000100101111100011011100111;
#4;
res_eth <= 32'b00010100101001010111001000010101;
#4;
res_eth <= 32'b00110111001000001110001100101001;
#4;
res_eth <= 32'b00011001010000101010000010100101;
#4;
res_eth <= 32'b00111011100011011000000001100011;
#4;
res_eth <= 32'b00011101111001110100111001010001;
#4;
res_eth <= 32'b00000010011010000011010111000010;
#4;
res_eth <= 32'b00100100100110100101001110101010;
#4;
res_eth <= 32'b01000111110110011100101110011011;
#4;
res_eth <= 32'b00101001110100100111110000110110;
#4;
res_eth <= 32'b00001101000010101000000001110010;
#4;
res_eth <= 32'b00101111110001110001101101010110;
#4;
res_eth <= 32'b01010010000011101011001010110001;
#4;
res_eth <= 32'b00110011101001100000001111010110;
#4;
res_eth <= 32'b00010111100110100100001010110000;
#4;
res_eth <= 32'b00111011011000101111011001011110;
#4;
res_eth <= 32'b01011101000011001011101000001001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01100001111111001000110111110101;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00100111110110111110110110011010;
#4;
res_eth <= 32'b01001011000101001001110010010001;
#4;
res_eth <= 32'b00101101100110010001100010000100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00110011101101111000111000011001;
#4;
res_eth <= 32'b00010110101111001111000101011100;
#4;
res_eth <= 32'b00111000110110011101010111010000;
#4;
res_eth <= 32'b01011011111001000101110110010010;
#4;
res_eth <= 32'b01111110001001100010100001100000;
#4;
res_eth <= 32'b00100001010001001000101000000000;
#4;
res_eth <= 32'b01000100001001101001000101010110;
#4;
res_eth <= 32'b01100101011111100110010101111111;
#4;
res_eth <= 32'b00001010001110001001100001111010;
#4;
res_eth <= 32'b01101010100101000101100001011011;
#4;
res_eth <= 32'b01001110101100100011011010110101;
#4;
res_eth <= 32'b01110000101011010101001111101000;
#4;
res_eth <= 32'b01010011111100001010110100101100;
#4;
res_eth <= 32'b00110110011100000001110111011010;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00000000000000000001010001001100;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01000000010111000001011010101100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00000111010100000011111001011001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00001011111111000000010110101100;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b01110101100011010001011110100011;
#4;
res_eth <= 32'b00011000001111010000100010011100;
#4;
res_eth <= 32'b01111001101010011011001101000111;
#4;
res_eth <= 32'b01011110010111001011001111010011;
#4;
res_eth <= 32'b01000000000010010111101110011000;
#4;
res_eth <= 32'b01100100010001000000101110000000;
#4;
res_eth <= 32'b00000101010100001110100001100101;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00001011010111100001000111000110;
#4;
res_eth <= 32'b00101101111100000110111010100011;
#4;
res_eth <= 32'b01001111000101101111011010001000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b00010101011101001011111011111100;
#4;
res_eth <= 32'b00000000000000000000000010001111;
#4;
res_eth <= 32'b01011011110010110100111010111010;
#4;
res_eth <= 32'b00111110001001001001101111100100;
#4;
res_eth <= 32'b00100001010010011110000001110001;
#4;
res_eth <= 32'b01111111100000000000000000000000;
#4;
res_eth <= 32'b00000000000000000000000000000000;
#4;
res_eth <= 32'b01001001100001001000011111000101;
#4;
res_eth <= 32'b01101100010001100011110011100011;
#4;
res_eth <= 32'b01001111111101011010110010000100;
#4;


end

reg [1:0]   opcode=0, rmode=0;
wire[31:0]  result;


always @(negedge clk) begin
    if(result != res_eth)
        $stop();
end
initial 
begin
    $dumpfile("out.vcd");
    $dumpvars(0, fmul_top);
    #1000000;
    $display ("SUCCESS");

    $finish();
end
endmodule
