`timescale 1ns/1ps


module testbench;
reg  [7:0] in;
wire [2:0] pow;

encoder #(.IN_SIZE(8)) DUT (
        .in(in),
        .pow(pow)
);

initial begin
$dumpfile("out.vcd");
$dumpvars(0,testbench);

	in = 8'b00000100;
	#10;

	in = 8'b00000010;
	#10;

	in = 8'b00010000;
	#10;

	in = 8'b10000000;
	#10;

$finish;
end
endmodule
